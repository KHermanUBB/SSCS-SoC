VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.470 3517.600 2030.030 3524.800 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3235.180 2924.800 3236.380 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1120.380 2924.800 1121.580 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.190 -4.800 2113.750 2.400 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.110 3517.600 2229.670 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 381.900 2924.800 383.100 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.190 -4.800 549.750 2.400 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.070 -4.800 332.630 2.400 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2728.670 -4.800 2729.230 2.400 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2842.140 2924.800 2843.340 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.790 3517.600 1796.350 3524.800 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 761.340 2.400 762.540 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 725.980 2924.800 727.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.030 3517.600 2046.590 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.390 3517.600 2628.950 3524.800 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.390 -4.800 1064.950 2.400 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.260 2924.800 3138.460 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3505.820 2924.800 3507.020 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.270 3517.600 65.830 3524.800 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.750 3517.600 1164.310 3524.800 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2631.340 2.400 2632.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 3517.600 1480.790 3524.800 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3099.180 2.400 3100.380 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2680.300 2.400 2681.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 455.340 2924.800 456.540 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 490.700 2.400 491.900 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2817.660 2924.800 2818.860 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2915.580 2924.800 2916.780 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 244.540 2.400 245.740 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1193.820 2924.800 1195.020 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.590 3517.600 2362.150 3524.800 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.110 3517.600 964.670 3524.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.230 3517.600 997.790 3524.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.430 3517.600 431.990 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 3517.600 98.950 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.510 3517.600 1098.070 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2755.100 2.400 2756.300 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.070 3517.600 1114.630 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.150 3517.600 331.710 3524.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.710 -4.800 1797.270 2.400 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2669.420 2924.800 2670.620 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 528.780 2924.800 529.980 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.030 -4.800 965.590 2.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.470 3517.600 1547.030 3524.800 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 86.780 2924.800 87.980 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 48.700 2.400 49.900 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2065.580 2.400 2066.780 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2844.590 3517.600 2845.150 3524.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 406.380 2924.800 407.580 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3296.380 2.400 3297.580 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2861.150 3517.600 2861.710 3524.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.070 3517.600 631.630 3524.800 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 701.500 2924.800 702.700 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 3517.600 215.790 3524.800 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2062.590 3517.600 2063.150 3524.800 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.990 3517.600 1230.550 3524.800 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 308.460 2924.800 309.660 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 3517.600 2562.710 3524.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3492.220 2.400 3493.420 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.150 -4.800 1780.710 2.400 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1819.420 2.400 1820.620 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3481.340 2924.800 3482.540 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.750 -4.800 2130.310 2.400 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.950 -4.800 2047.510 2.400 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2778.350 3517.600 2778.910 3524.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.550 -4.800 649.110 2.400 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.590 -4.800 499.150 2.400 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2645.870 -4.800 2646.430 2.400 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1464.460 2924.800 1465.660 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2744.220 2924.800 2745.420 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2730.620 2.400 2731.820 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.470 -4.800 2214.030 2.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.950 -4.800 2829.510 2.400 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 3517.600 481.670 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.750 3517.600 2728.310 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 3517.600 16.150 3524.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 122.140 2.400 123.340 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.270 -4.800 1514.830 2.400 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 -4.800 83.310 2.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1672.540 2.400 1673.740 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2571.500 2924.800 2572.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1229.180 2.400 1230.380 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1316.220 2924.800 1317.420 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.750 3517.600 681.310 3524.800 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1031.980 2.400 1033.180 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2901.980 2.400 2903.180 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 3517.600 165.190 3524.800 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3112.780 2924.800 3113.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.510 3517.600 2662.070 3524.800 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 184.700 2924.800 185.900 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.270 3517.600 1629.830 3524.800 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.030 3517.600 781.590 3524.800 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.070 -4.800 1298.630 2.400 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3518.060 2.400 3519.260 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 3517.600 398.870 3524.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2866.620 2924.800 2867.820 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.510 3517.600 2179.070 3524.800 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2828.540 2.400 2829.740 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.710 -4.800 233.270 2.400 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.670 3517.600 1464.230 3524.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.990 -4.800 2380.550 2.400 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 541.020 2.400 542.220 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2557.900 2.400 2559.100 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.350 3517.600 248.910 3524.800 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2398.780 2924.800 2399.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.070 3517.600 2379.630 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 -4.800 249.830 2.400 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2287.260 2.400 2288.460 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1253.660 2.400 1254.860 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1686.140 2924.800 1687.340 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2311.740 2.400 2312.940 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.230 -4.800 399.790 2.400 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.670 3517.600 498.230 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.300 2924.800 2375.500 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.430 3517.600 1213.990 3524.800 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.150 3517.600 1596.710 3524.800 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.670 -4.800 1947.230 2.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.910 3517.600 1047.470 3524.800 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 357.420 2924.800 358.620 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2300.860 2924.800 2302.060 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.630 -4.800 349.190 2.400 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.830 -4.800 1048.390 2.400 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2227.420 2924.800 2228.620 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1415.500 2924.800 1416.700 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.430 -4.800 1880.990 2.400 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.790 -4.800 416.350 2.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2412.190 3517.600 2412.750 3524.800 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.670 -4.800 682.230 2.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.110 -4.800 665.670 2.400 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 -4.800 166.110 2.400 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2128.830 3517.600 2129.390 3524.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1180.220 2.400 1181.420 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2103.660 2924.800 2104.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.750 -4.800 1348.310 2.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 898.700 2924.800 899.900 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.940 2.400 2510.140 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.470 3517.600 1064.030 3524.800 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.510 3517.600 1397.070 3524.800 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.350 3517.600 1030.910 3524.800 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3285.500 2924.800 3286.700 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1242.780 2924.800 1243.980 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1106.780 2.400 1107.980 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 3517.600 265.470 3524.800 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1918.700 2.400 1919.900 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3247.420 2.400 3248.620 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.670 3517.600 981.230 3524.800 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 3517.600 365.750 3524.800 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.230 3517.600 1779.790 3524.800 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 195.580 2.400 196.780 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.470 -4.800 466.030 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2655.820 2.400 2657.020 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.910 -4.800 1714.470 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3334.460 2924.800 3335.660 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1340.700 2924.800 1341.900 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.390 -4.800 1547.950 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2202.940 2924.800 2204.140 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2139.020 2.400 2140.220 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.830 3517.600 1347.390 3524.800 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2522.540 2924.800 2523.740 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 3517.600 1263.670 3524.800 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2128.140 2924.800 2129.340 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1218.300 2924.800 1219.500 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.550 -4.800 1914.110 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 3517.600 2262.790 3524.800 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 62.300 2924.800 63.500 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1524.300 2.400 1525.500 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2251.900 2924.800 2253.100 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.670 3517.600 2545.230 3524.800 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.870 3517.600 1197.430 3524.800 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2644.940 2924.800 2646.140 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2712.110 -4.800 2712.670 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.990 -4.800 2679.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 3517.600 1763.230 3524.800 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3271.900 2.400 3273.100 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 811.660 2.400 812.860 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 111.260 2924.800 112.460 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2336.220 2.400 2337.420 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.750 3517.600 382.310 3524.800 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1426.380 2.400 1427.580 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 343.820 2.400 345.020 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 3517.600 1297.710 3524.800 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.670 -4.800 1165.230 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1562.380 2924.800 1563.580 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.150 3517.600 814.710 3524.800 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1131.260 2.400 1132.460 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 712.380 2.400 713.580 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.150 -4.800 998.710 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.710 3517.600 1613.270 3524.800 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3172.620 2.400 3173.820 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2926.460 2.400 2927.660 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 799.420 2924.800 800.620 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.870 -4.800 2163.430 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.910 -4.800 1231.470 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.550 3517.600 465.110 3524.800 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 3517.600 182.670 3524.800 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1637.180 2924.800 1638.380 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.710 3517.600 1314.270 3524.800 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.390 3517.600 880.950 3524.800 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 947.660 2924.800 948.860 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 319.340 2.400 320.540 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1808.540 2924.800 1809.740 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.100 2.400 1328.300 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1932.300 2924.800 1933.500 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2114.540 2.400 2115.740 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.630 3517.600 648.190 3524.800 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1730.470 -4.800 1731.030 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2877.710 3517.600 2878.270 3524.800 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2533.420 2.400 2534.620 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 3517.600 199.230 3524.800 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 417.260 2.400 418.460 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 -4.800 17.070 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2178.460 2924.800 2179.660 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2853.020 2.400 2854.220 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3088.300 2924.800 3089.500 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.110 -4.800 366.670 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1784.060 2924.800 1785.260 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.070 3517.600 1896.630 3524.800 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2079.180 2924.800 2080.380 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2545.590 -4.800 2546.150 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1611.340 2924.800 1612.540 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.870 3517.600 1979.430 3524.800 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2582.380 2.400 2583.580 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 3517.600 2762.350 3524.800 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2090.060 2.400 2091.260 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2976.780 2.400 2977.980 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.030 -4.800 2529.590 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 874.220 2924.800 875.420 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2768.700 2924.800 2769.900 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2990.380 2924.800 2991.580 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.350 3517.600 2295.910 3524.800 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 392.780 2.400 393.980 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1021.100 2924.800 1022.300 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 37.820 2924.800 39.020 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2528.110 3517.600 2528.670 3524.800 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.550 -4.800 1431.110 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2693.900 2924.800 2695.100 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 466.220 2.400 467.420 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2629.310 -4.800 2629.870 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1144.860 2924.800 1146.060 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.070 3517.600 2678.630 3524.800 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.950 -4.800 2346.510 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.310 3517.600 1180.870 3524.800 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1759.580 2924.800 1760.780 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2245.670 3517.600 2246.230 3524.800 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.030 3517.600 1080.590 3524.800 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.630 3517.600 1913.190 3524.800 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1992.140 2.400 1993.340 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2296.270 -4.800 2296.830 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2262.780 2.400 2263.980 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2595.980 2924.800 2597.180 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 3517.600 1430.190 3524.800 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1745.980 2.400 1747.180 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3186.220 2924.800 3187.420 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2804.060 2.400 2805.260 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.270 3517.600 2112.830 3524.800 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.110 -4.800 1148.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3050.220 2.400 3051.420 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1513.420 2924.800 1514.620 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.950 3517.600 1863.510 3524.800 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1881.980 2924.800 1883.180 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.150 -4.800 515.710 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 652.540 2924.800 653.740 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.270 3517.600 2595.830 3524.800 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 283.980 2924.800 285.180 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.990 -4.800 632.550 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1439.980 2924.800 1441.180 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2152.620 2924.800 2153.820 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.550 3517.600 2213.110 3524.800 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.270 -4.800 1813.830 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1648.060 2.400 1649.260 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 504.300 2924.800 505.500 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.630 -4.800 832.190 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.990 3517.600 448.550 3524.800 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 258.140 2924.800 259.340 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.790 -4.800 1681.350 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.790 3517.600 531.350 3524.800 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1488.940 2924.800 1490.140 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2495.910 -4.800 2496.470 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 825.260 2924.800 826.460 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 885.100 2.400 886.300 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.950 -4.800 1081.510 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 171.100 2.400 172.300 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3161.740 2924.800 3162.940 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2711.190 3517.600 2711.750 3524.800 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 3517.600 298.590 3524.800 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.470 3517.600 765.030 3524.800 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.310 3517.600 697.870 3524.800 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.910 -4.800 932.470 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.070 -4.800 2563.630 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 3517.600 82.390 3524.800 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2779.580 2.400 2780.780 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1981.260 2924.800 1982.460 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1710.620 2924.800 1711.820 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1082.300 2.400 1083.500 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.350 3517.600 731.910 3524.800 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2762.710 -4.800 2763.270 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.430 3517.600 1696.990 3524.800 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 554.620 2924.800 555.820 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3197.100 2.400 3198.300 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 579.100 2924.800 580.300 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2462.790 -4.800 2463.350 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.830 3517.600 2612.390 3524.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2238.300 2.400 2239.500 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.710 3517.600 831.270 3524.800 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.510 -4.800 1282.070 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.030 -4.800 1264.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.790 -4.800 1980.350 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 3517.600 1663.870 3524.800 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1450.860 2.400 1452.060 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1770.460 2.400 1771.660 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.190 3517.600 1929.750 3524.800 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 135.740 2924.800 136.940 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.190 3517.600 664.750 3524.800 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.230 -4.800 2446.790 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2695.550 -4.800 2696.110 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 13.340 2924.800 14.540 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.550 3517.600 1247.110 3524.800 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1267.260 2924.800 1268.460 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 565.500 2.400 566.700 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 3517.600 348.270 3524.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 368.300 2.400 369.500 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1967.660 2.400 1968.860 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.950 -4.800 1564.510 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.950 3517.600 897.510 3524.800 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 -4.800 282.950 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.870 3517.600 1680.430 3524.800 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 3517.600 232.350 3524.800 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 3517.600 2645.510 3524.800 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1475.340 2.400 1476.540 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 515.180 2.400 516.380 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 3517.600 2096.270 3524.800 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2435.500 2.400 2436.700 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.190 -4.800 848.750 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.030 -4.800 1747.590 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.590 3517.600 1281.150 3524.800 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.510 3517.600 615.070 3524.800 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1943.180 2.400 1944.380 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.150 -4.800 1481.710 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.110 -4.800 1447.670 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.550 3517.600 2512.110 3524.800 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 736.860 2.400 738.060 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.750 3517.600 2429.310 3524.800 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2484.460 2.400 2485.660 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.430 -4.800 2179.990 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2429.670 -4.800 2430.230 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1956.780 2924.800 1957.980 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 677.020 2924.800 678.220 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.830 3517.600 864.390 3524.800 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.190 -4.800 1331.750 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.230 -4.800 1963.790 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.710 -4.800 1015.270 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 3517.600 115.510 3524.800 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.710 -4.800 1498.270 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.070 -4.800 2080.630 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.230 -4.800 1664.790 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.270 -4.800 732.830 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.390 3517.600 581.950 3524.800 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.870 -4.800 1381.430 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 614.460 2.400 615.660 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2612.750 -4.800 2613.310 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 628.060 2924.800 629.260 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.430 3517.600 914.990 3524.800 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 294.860 2.400 296.060 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3418.780 2.400 3419.980 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1302.620 2.400 1303.820 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 3517.600 2745.790 3524.800 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.590 -4.800 2247.150 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3407.900 2924.800 3409.100 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 687.900 2.400 689.100 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2746.150 -4.800 2746.710 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1857.500 2924.800 1858.700 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3320.860 2.400 3322.060 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.630 3517.600 1131.190 3524.800 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.190 3517.600 1446.750 3524.800 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510 3517.600 132.070 3524.800 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.510 -4.800 2064.070 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.390 -4.800 2329.950 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.590 3517.600 1580.150 3524.800 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.510 -4.800 799.070 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2894.270 3517.600 2894.830 3524.800 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1868.380 2.400 1869.580 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1697.020 2.400 1698.220 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.030 3517.600 2345.590 3524.800 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.790 3517.600 2279.350 3524.800 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.270 -4.800 2779.830 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.470 -4.800 1248.030 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.470 3517.600 282.030 3524.800 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2811.470 3517.600 2812.030 3524.800 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 233.660 2924.800 234.860 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.470 3517.600 2329.030 3524.800 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.790 -4.800 715.350 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 909.580 2.400 910.780 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.830 -4.800 2014.390 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2694.630 3517.600 2695.190 3524.800 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3074.700 2.400 3075.900 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3467.740 2.400 3468.940 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.950 3517.600 2162.510 3524.800 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.430 -4.800 1098.990 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2793.180 2924.800 2794.380 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.350 -4.800 1996.910 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1833.020 2924.800 1834.220 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.750 3517.600 1647.310 3524.800 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.070 -4.800 1597.630 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.990 -4.800 1414.550 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1721.500 2.400 1722.700 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1291.740 2924.800 1292.940 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.870 3517.600 415.430 3524.800 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2005.740 2924.800 2006.940 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.910 3517.600 748.470 3524.800 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.590 -4.800 982.150 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 3517.600 1746.670 3524.800 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1352.940 2.400 1354.140 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1070.060 2924.800 1071.260 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1661.660 2924.800 1662.860 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.150 -4.800 2263.710 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 750.460 2924.800 751.660 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2473.580 2924.800 2474.780 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.550 3517.600 1730.110 3524.800 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 934.060 2.400 935.260 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 441.740 2.400 442.940 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.950 -4.800 782.510 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.860 2924.800 432.060 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 -4.800 183.590 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.070 -4.800 815.630 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 332.940 2924.800 334.140 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3432.380 2924.800 3433.580 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1391.020 2924.800 1392.220 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.950 -4.800 299.510 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1095.900 2924.800 1097.100 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.990 -4.800 1897.550 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.870 3517.600 2462.430 3524.800 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.590 -4.800 1764.150 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1907.820 2924.800 1909.020 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2794.910 3517.600 2795.470 3524.800 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1401.900 2.400 1403.100 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3001.260 2.400 3002.460 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 3517.600 2828.590 3524.800 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 589.980 2.400 591.180 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1843.900 2.400 1845.100 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2911.750 -4.800 2912.310 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1155.740 2.400 1156.940 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1573.260 2.400 1574.460 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.070 3517.600 1413.630 3524.800 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.630 -4.800 2097.190 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2385.180 2.400 2386.380 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2041.100 2.400 2042.300 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2016.620 2.400 2017.820 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3309.980 2924.800 3311.180 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.470 -4.800 2513.030 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 983.020 2.400 984.220 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.110 -4.800 2413.670 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 958.540 2.400 959.740 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.030 -4.800 482.590 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.830 -4.800 749.390 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.190 -4.800 2596.750 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 923.180 2924.800 924.380 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2964.540 2924.800 2965.740 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.790 3517.600 1497.350 3524.800 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 3517.600 1380.510 3524.800 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2950.940 2.400 2952.140 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.350 -4.800 915.910 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3358.940 2924.800 3360.140 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1794.940 2.400 1796.140 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.590 3517.600 798.150 3524.800 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.310 -4.800 582.870 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2891.100 2924.800 2892.300 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 785.820 2.400 787.020 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.830 3517.600 1830.390 3524.800 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.910 3517.600 2312.470 3524.800 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.310 3517.600 2445.870 3524.800 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2478.430 3517.600 2478.990 3524.800 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 270.380 2.400 271.580 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 3517.600 1563.590 3524.800 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 -4.800 99.870 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.070 -4.800 33.630 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 638.940 2.400 640.140 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 479.820 2924.800 481.020 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2706.140 2.400 2707.340 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2606.860 2.400 2608.060 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3148.140 2.400 3149.340 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1623.580 2.400 1624.780 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1377.420 2.400 1378.620 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1056.460 2.400 1057.660 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.350 3517.600 1513.910 3524.800 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.230 -4.800 1181.790 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3025.740 2.400 3026.940 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2449.100 2924.800 2450.300 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3261.020 2924.800 3262.220 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 146.620 2.400 147.820 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 160.220 2924.800 161.420 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3063.820 2924.800 3065.020 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.190 3517.600 1147.750 3524.800 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2498.060 2924.800 2499.260 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.830 -4.800 2313.390 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.350 3517.600 1812.910 3524.800 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 603.580 2924.800 604.780 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.550 3517.600 948.110 3524.800 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2795.830 -4.800 2796.390 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3394.300 2.400 3395.500 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.670 -4.800 383.230 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2349.820 2924.800 2351.020 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3014.860 2924.800 3016.060 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.390 -4.800 765.950 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 3517.600 148.630 3524.800 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1894.220 2.400 1895.420 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 860.620 2.400 861.820 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 3517.600 49.270 3524.800 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 3517.600 315.150 3524.800 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3369.820 2.400 3371.020 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1586.860 2924.800 1588.060 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.270 3517.600 1330.830 3524.800 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.870 3517.600 714.430 3524.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2877.500 2.400 2878.700 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 -4.800 266.390 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2213.820 2.400 2215.020 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3210.700 2924.800 3211.900 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2940.060 2924.800 2941.260 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2620.460 2924.800 2621.660 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1366.540 2924.800 1367.740 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2812.390 -4.800 2812.950 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.390 3517.600 1363.950 3524.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1278.140 2.400 1279.340 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.670 -4.800 1648.230 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.510 -4.800 2363.070 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 972.140 2924.800 973.340 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3345.340 2.400 3346.540 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.510 -4.800 1581.070 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.510 -4.800 316.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.270 3517.600 548.830 3524.800 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2423.260 2924.800 2424.460 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2578.710 3517.600 2579.270 3524.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.990 -4.800 1115.550 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.510 3517.600 1880.070 3524.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1735.100 2924.800 1736.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.030 -4.800 2230.590 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.390 3517.600 1846.950 3524.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 663.420 2.400 664.620 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.870 -4.800 898.430 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.990 -4.800 149.550 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.070 -4.800 2862.630 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1045.580 2924.800 1046.780 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.950 3517.600 598.510 3524.800 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 3517.600 2911.390 3524.800 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2164.860 2.400 2166.060 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2459.980 2.400 2461.180 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2360.700 2.400 2361.900 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 -4.800 116.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.430 -4.800 615.990 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2030.220 2924.800 2031.420 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 220.060 2.400 221.260 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.990 3517.600 1713.550 3524.800 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.630 3517.600 2396.190 3524.800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3443.260 2.400 3444.460 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.350 -4.800 432.910 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2325.340 2924.800 2326.540 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.990 3517.600 2495.550 3524.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1597.740 2.400 1598.940 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3039.340 2924.800 3040.540 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1169.340 2924.800 1170.540 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 97.660 2.400 98.860 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.990 3517.600 2196.550 3524.800 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.830 3517.600 565.390 3524.800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.310 -4.800 881.870 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2276.380 2924.800 2277.580 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.710 -4.800 2280.270 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 996.620 2924.800 997.820 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1499.820 2.400 1501.020 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2878.630 -4.800 2879.190 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.910 -4.800 449.470 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 24.220 2.400 25.420 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.390 3517.600 2145.950 3524.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3383.420 2924.800 3384.620 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2895.190 -4.800 2895.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 -4.800 216.710 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2054.700 2924.800 2055.900 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 -4.800 66.750 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3456.860 2924.800 3458.060 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2079.150 3517.600 2079.710 3524.800 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 209.180 2924.800 210.380 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.430 3517.600 1995.990 3524.800 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.310 -4.800 1847.870 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 73.180 2.400 74.380 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.750 -4.800 1831.310 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 -4.800 0.510 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.310 -4.800 2146.870 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1548.780 2.400 1549.980 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.270 3517.600 847.830 3524.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1007.500 2.400 1008.700 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.750 -4.800 566.310 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 -4.800 200.150 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.910 3517.600 1530.470 3524.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.990 3517.600 931.550 3524.800 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.590 -4.800 1465.150 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.910 3517.600 2013.470 3524.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 774.940 2924.800 776.140 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2409.660 2.400 2410.860 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2719.740 2924.800 2720.940 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.870 -4.800 599.430 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.630 -4.800 1614.190 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2547.020 2924.800 2548.220 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.190 -4.800 1630.750 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.310 3517.600 1962.870 3524.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.750 3517.600 1946.310 3524.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 3517.600 32.710 3524.800 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.230 3517.600 514.790 3524.800 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.110 -4.800 1930.670 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 836.140 2.400 837.340 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3221.580 2.400 3222.780 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1537.900 2924.800 1539.100 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 194.725 14.025 2723.515 3320.355 ;
      LAYER met1 ;
        RECT 0.070 13.980 2912.190 3515.220 ;
      LAYER met2 ;
        RECT 0.100 3517.320 15.310 3518.845 ;
        RECT 16.430 3517.320 31.870 3518.845 ;
        RECT 32.990 3517.320 48.430 3518.845 ;
        RECT 49.550 3517.320 64.990 3518.845 ;
        RECT 66.110 3517.320 81.550 3518.845 ;
        RECT 82.670 3517.320 98.110 3518.845 ;
        RECT 99.230 3517.320 114.670 3518.845 ;
        RECT 115.790 3517.320 131.230 3518.845 ;
        RECT 132.350 3517.320 147.790 3518.845 ;
        RECT 148.910 3517.320 164.350 3518.845 ;
        RECT 165.470 3517.320 181.830 3518.845 ;
        RECT 182.950 3517.320 198.390 3518.845 ;
        RECT 199.510 3517.320 214.950 3518.845 ;
        RECT 216.070 3517.320 231.510 3518.845 ;
        RECT 232.630 3517.320 248.070 3518.845 ;
        RECT 249.190 3517.320 264.630 3518.845 ;
        RECT 265.750 3517.320 281.190 3518.845 ;
        RECT 282.310 3517.320 297.750 3518.845 ;
        RECT 298.870 3517.320 314.310 3518.845 ;
        RECT 315.430 3517.320 330.870 3518.845 ;
        RECT 331.990 3517.320 347.430 3518.845 ;
        RECT 348.550 3517.320 364.910 3518.845 ;
        RECT 366.030 3517.320 381.470 3518.845 ;
        RECT 382.590 3517.320 398.030 3518.845 ;
        RECT 399.150 3517.320 414.590 3518.845 ;
        RECT 415.710 3517.320 431.150 3518.845 ;
        RECT 432.270 3517.320 447.710 3518.845 ;
        RECT 448.830 3517.320 464.270 3518.845 ;
        RECT 465.390 3517.320 480.830 3518.845 ;
        RECT 481.950 3517.320 497.390 3518.845 ;
        RECT 498.510 3517.320 513.950 3518.845 ;
        RECT 515.070 3517.320 530.510 3518.845 ;
        RECT 531.630 3517.320 547.990 3518.845 ;
        RECT 549.110 3517.320 564.550 3518.845 ;
        RECT 565.670 3517.320 581.110 3518.845 ;
        RECT 582.230 3517.320 597.670 3518.845 ;
        RECT 598.790 3517.320 614.230 3518.845 ;
        RECT 615.350 3517.320 630.790 3518.845 ;
        RECT 631.910 3517.320 647.350 3518.845 ;
        RECT 648.470 3517.320 663.910 3518.845 ;
        RECT 665.030 3517.320 680.470 3518.845 ;
        RECT 681.590 3517.320 697.030 3518.845 ;
        RECT 698.150 3517.320 713.590 3518.845 ;
        RECT 714.710 3517.320 731.070 3518.845 ;
        RECT 732.190 3517.320 747.630 3518.845 ;
        RECT 748.750 3517.320 764.190 3518.845 ;
        RECT 765.310 3517.320 780.750 3518.845 ;
        RECT 781.870 3517.320 797.310 3518.845 ;
        RECT 798.430 3517.320 813.870 3518.845 ;
        RECT 814.990 3517.320 830.430 3518.845 ;
        RECT 831.550 3517.320 846.990 3518.845 ;
        RECT 848.110 3517.320 863.550 3518.845 ;
        RECT 864.670 3517.320 880.110 3518.845 ;
        RECT 881.230 3517.320 896.670 3518.845 ;
        RECT 897.790 3517.320 914.150 3518.845 ;
        RECT 915.270 3517.320 930.710 3518.845 ;
        RECT 931.830 3517.320 947.270 3518.845 ;
        RECT 948.390 3517.320 963.830 3518.845 ;
        RECT 964.950 3517.320 980.390 3518.845 ;
        RECT 981.510 3517.320 996.950 3518.845 ;
        RECT 998.070 3517.320 1013.510 3518.845 ;
        RECT 1014.630 3517.320 1030.070 3518.845 ;
        RECT 1031.190 3517.320 1046.630 3518.845 ;
        RECT 1047.750 3517.320 1063.190 3518.845 ;
        RECT 1064.310 3517.320 1079.750 3518.845 ;
        RECT 1080.870 3517.320 1097.230 3518.845 ;
        RECT 1098.350 3517.320 1113.790 3518.845 ;
        RECT 1114.910 3517.320 1130.350 3518.845 ;
        RECT 1131.470 3517.320 1146.910 3518.845 ;
        RECT 1148.030 3517.320 1163.470 3518.845 ;
        RECT 1164.590 3517.320 1180.030 3518.845 ;
        RECT 1181.150 3517.320 1196.590 3518.845 ;
        RECT 1197.710 3517.320 1213.150 3518.845 ;
        RECT 1214.270 3517.320 1229.710 3518.845 ;
        RECT 1230.830 3517.320 1246.270 3518.845 ;
        RECT 1247.390 3517.320 1262.830 3518.845 ;
        RECT 1263.950 3517.320 1280.310 3518.845 ;
        RECT 1281.430 3517.320 1296.870 3518.845 ;
        RECT 1297.990 3517.320 1313.430 3518.845 ;
        RECT 1314.550 3517.320 1329.990 3518.845 ;
        RECT 1331.110 3517.320 1346.550 3518.845 ;
        RECT 1347.670 3517.320 1363.110 3518.845 ;
        RECT 1364.230 3517.320 1379.670 3518.845 ;
        RECT 1380.790 3517.320 1396.230 3518.845 ;
        RECT 1397.350 3517.320 1412.790 3518.845 ;
        RECT 1413.910 3517.320 1429.350 3518.845 ;
        RECT 1430.470 3517.320 1445.910 3518.845 ;
        RECT 1447.030 3517.320 1463.390 3518.845 ;
        RECT 1464.510 3517.320 1479.950 3518.845 ;
        RECT 1481.070 3517.320 1496.510 3518.845 ;
        RECT 1497.630 3517.320 1513.070 3518.845 ;
        RECT 1514.190 3517.320 1529.630 3518.845 ;
        RECT 1530.750 3517.320 1546.190 3518.845 ;
        RECT 1547.310 3517.320 1562.750 3518.845 ;
        RECT 1563.870 3517.320 1579.310 3518.845 ;
        RECT 1580.430 3517.320 1595.870 3518.845 ;
        RECT 1596.990 3517.320 1612.430 3518.845 ;
        RECT 1613.550 3517.320 1628.990 3518.845 ;
        RECT 1630.110 3517.320 1646.470 3518.845 ;
        RECT 1647.590 3517.320 1663.030 3518.845 ;
        RECT 1664.150 3517.320 1679.590 3518.845 ;
        RECT 1680.710 3517.320 1696.150 3518.845 ;
        RECT 1697.270 3517.320 1712.710 3518.845 ;
        RECT 1713.830 3517.320 1729.270 3518.845 ;
        RECT 1730.390 3517.320 1745.830 3518.845 ;
        RECT 1746.950 3517.320 1762.390 3518.845 ;
        RECT 1763.510 3517.320 1778.950 3518.845 ;
        RECT 1780.070 3517.320 1795.510 3518.845 ;
        RECT 1796.630 3517.320 1812.070 3518.845 ;
        RECT 1813.190 3517.320 1829.550 3518.845 ;
        RECT 1830.670 3517.320 1846.110 3518.845 ;
        RECT 1847.230 3517.320 1862.670 3518.845 ;
        RECT 1863.790 3517.320 1879.230 3518.845 ;
        RECT 1880.350 3517.320 1895.790 3518.845 ;
        RECT 1896.910 3517.320 1912.350 3518.845 ;
        RECT 1913.470 3517.320 1928.910 3518.845 ;
        RECT 1930.030 3517.320 1945.470 3518.845 ;
        RECT 1946.590 3517.320 1962.030 3518.845 ;
        RECT 1963.150 3517.320 1978.590 3518.845 ;
        RECT 1979.710 3517.320 1995.150 3518.845 ;
        RECT 1996.270 3517.320 2012.630 3518.845 ;
        RECT 2013.750 3517.320 2029.190 3518.845 ;
        RECT 2030.310 3517.320 2045.750 3518.845 ;
        RECT 2046.870 3517.320 2062.310 3518.845 ;
        RECT 2063.430 3517.320 2078.870 3518.845 ;
        RECT 2079.990 3517.320 2095.430 3518.845 ;
        RECT 2096.550 3517.320 2111.990 3518.845 ;
        RECT 2113.110 3517.320 2128.550 3518.845 ;
        RECT 2129.670 3517.320 2145.110 3518.845 ;
        RECT 2146.230 3517.320 2161.670 3518.845 ;
        RECT 2162.790 3517.320 2178.230 3518.845 ;
        RECT 2179.350 3517.320 2195.710 3518.845 ;
        RECT 2196.830 3517.320 2212.270 3518.845 ;
        RECT 2213.390 3517.320 2228.830 3518.845 ;
        RECT 2229.950 3517.320 2245.390 3518.845 ;
        RECT 2246.510 3517.320 2261.950 3518.845 ;
        RECT 2263.070 3517.320 2278.510 3518.845 ;
        RECT 2279.630 3517.320 2295.070 3518.845 ;
        RECT 2296.190 3517.320 2311.630 3518.845 ;
        RECT 2312.750 3517.320 2328.190 3518.845 ;
        RECT 2329.310 3517.320 2344.750 3518.845 ;
        RECT 2345.870 3517.320 2361.310 3518.845 ;
        RECT 2362.430 3517.320 2378.790 3518.845 ;
        RECT 2379.910 3517.320 2395.350 3518.845 ;
        RECT 2396.470 3517.320 2411.910 3518.845 ;
        RECT 2413.030 3517.320 2428.470 3518.845 ;
        RECT 2429.590 3517.320 2445.030 3518.845 ;
        RECT 2446.150 3517.320 2461.590 3518.845 ;
        RECT 2462.710 3517.320 2478.150 3518.845 ;
        RECT 2479.270 3517.320 2494.710 3518.845 ;
        RECT 2495.830 3517.320 2511.270 3518.845 ;
        RECT 2512.390 3517.320 2527.830 3518.845 ;
        RECT 2528.950 3517.320 2544.390 3518.845 ;
        RECT 2545.510 3517.320 2561.870 3518.845 ;
        RECT 2562.990 3517.320 2578.430 3518.845 ;
        RECT 2579.550 3517.320 2594.990 3518.845 ;
        RECT 2596.110 3517.320 2611.550 3518.845 ;
        RECT 2612.670 3517.320 2628.110 3518.845 ;
        RECT 2629.230 3517.320 2644.670 3518.845 ;
        RECT 2645.790 3517.320 2661.230 3518.845 ;
        RECT 2662.350 3517.320 2677.790 3518.845 ;
        RECT 2678.910 3517.320 2694.350 3518.845 ;
        RECT 2695.470 3517.320 2710.910 3518.845 ;
        RECT 2712.030 3517.320 2727.470 3518.845 ;
        RECT 2728.590 3517.320 2744.950 3518.845 ;
        RECT 2746.070 3517.320 2761.510 3518.845 ;
        RECT 2762.630 3517.320 2778.070 3518.845 ;
        RECT 2779.190 3517.320 2794.630 3518.845 ;
        RECT 2795.750 3517.320 2811.190 3518.845 ;
        RECT 2812.310 3517.320 2827.750 3518.845 ;
        RECT 2828.870 3517.320 2844.310 3518.845 ;
        RECT 2845.430 3517.320 2860.870 3518.845 ;
        RECT 2861.990 3517.320 2877.430 3518.845 ;
        RECT 2878.550 3517.320 2893.990 3518.845 ;
        RECT 2895.110 3517.320 2910.550 3518.845 ;
        RECT 2911.670 3517.320 2912.160 3518.845 ;
        RECT 0.100 2.680 2912.160 3517.320 ;
        RECT 0.790 2.310 16.230 2.680 ;
        RECT 17.350 2.310 32.790 2.680 ;
        RECT 33.910 2.310 49.350 2.680 ;
        RECT 50.470 2.310 65.910 2.680 ;
        RECT 67.030 2.310 82.470 2.680 ;
        RECT 83.590 2.310 99.030 2.680 ;
        RECT 100.150 2.310 115.590 2.680 ;
        RECT 116.710 2.310 132.150 2.680 ;
        RECT 133.270 2.310 148.710 2.680 ;
        RECT 149.830 2.310 165.270 2.680 ;
        RECT 166.390 2.310 182.750 2.680 ;
        RECT 183.870 2.310 199.310 2.680 ;
        RECT 200.430 2.310 215.870 2.680 ;
        RECT 216.990 2.310 232.430 2.680 ;
        RECT 233.550 2.310 248.990 2.680 ;
        RECT 250.110 2.310 265.550 2.680 ;
        RECT 266.670 2.310 282.110 2.680 ;
        RECT 283.230 2.310 298.670 2.680 ;
        RECT 299.790 2.310 315.230 2.680 ;
        RECT 316.350 2.310 331.790 2.680 ;
        RECT 332.910 2.310 348.350 2.680 ;
        RECT 349.470 2.310 365.830 2.680 ;
        RECT 366.950 2.310 382.390 2.680 ;
        RECT 383.510 2.310 398.950 2.680 ;
        RECT 400.070 2.310 415.510 2.680 ;
        RECT 416.630 2.310 432.070 2.680 ;
        RECT 433.190 2.310 448.630 2.680 ;
        RECT 449.750 2.310 465.190 2.680 ;
        RECT 466.310 2.310 481.750 2.680 ;
        RECT 482.870 2.310 498.310 2.680 ;
        RECT 499.430 2.310 514.870 2.680 ;
        RECT 515.990 2.310 531.430 2.680 ;
        RECT 532.550 2.310 548.910 2.680 ;
        RECT 550.030 2.310 565.470 2.680 ;
        RECT 566.590 2.310 582.030 2.680 ;
        RECT 583.150 2.310 598.590 2.680 ;
        RECT 599.710 2.310 615.150 2.680 ;
        RECT 616.270 2.310 631.710 2.680 ;
        RECT 632.830 2.310 648.270 2.680 ;
        RECT 649.390 2.310 664.830 2.680 ;
        RECT 665.950 2.310 681.390 2.680 ;
        RECT 682.510 2.310 697.950 2.680 ;
        RECT 699.070 2.310 714.510 2.680 ;
        RECT 715.630 2.310 731.990 2.680 ;
        RECT 733.110 2.310 748.550 2.680 ;
        RECT 749.670 2.310 765.110 2.680 ;
        RECT 766.230 2.310 781.670 2.680 ;
        RECT 782.790 2.310 798.230 2.680 ;
        RECT 799.350 2.310 814.790 2.680 ;
        RECT 815.910 2.310 831.350 2.680 ;
        RECT 832.470 2.310 847.910 2.680 ;
        RECT 849.030 2.310 864.470 2.680 ;
        RECT 865.590 2.310 881.030 2.680 ;
        RECT 882.150 2.310 897.590 2.680 ;
        RECT 898.710 2.310 915.070 2.680 ;
        RECT 916.190 2.310 931.630 2.680 ;
        RECT 932.750 2.310 948.190 2.680 ;
        RECT 949.310 2.310 964.750 2.680 ;
        RECT 965.870 2.310 981.310 2.680 ;
        RECT 982.430 2.310 997.870 2.680 ;
        RECT 998.990 2.310 1014.430 2.680 ;
        RECT 1015.550 2.310 1030.990 2.680 ;
        RECT 1032.110 2.310 1047.550 2.680 ;
        RECT 1048.670 2.310 1064.110 2.680 ;
        RECT 1065.230 2.310 1080.670 2.680 ;
        RECT 1081.790 2.310 1098.150 2.680 ;
        RECT 1099.270 2.310 1114.710 2.680 ;
        RECT 1115.830 2.310 1131.270 2.680 ;
        RECT 1132.390 2.310 1147.830 2.680 ;
        RECT 1148.950 2.310 1164.390 2.680 ;
        RECT 1165.510 2.310 1180.950 2.680 ;
        RECT 1182.070 2.310 1197.510 2.680 ;
        RECT 1198.630 2.310 1214.070 2.680 ;
        RECT 1215.190 2.310 1230.630 2.680 ;
        RECT 1231.750 2.310 1247.190 2.680 ;
        RECT 1248.310 2.310 1263.750 2.680 ;
        RECT 1264.870 2.310 1281.230 2.680 ;
        RECT 1282.350 2.310 1297.790 2.680 ;
        RECT 1298.910 2.310 1314.350 2.680 ;
        RECT 1315.470 2.310 1330.910 2.680 ;
        RECT 1332.030 2.310 1347.470 2.680 ;
        RECT 1348.590 2.310 1364.030 2.680 ;
        RECT 1365.150 2.310 1380.590 2.680 ;
        RECT 1381.710 2.310 1397.150 2.680 ;
        RECT 1398.270 2.310 1413.710 2.680 ;
        RECT 1414.830 2.310 1430.270 2.680 ;
        RECT 1431.390 2.310 1446.830 2.680 ;
        RECT 1447.950 2.310 1464.310 2.680 ;
        RECT 1465.430 2.310 1480.870 2.680 ;
        RECT 1481.990 2.310 1497.430 2.680 ;
        RECT 1498.550 2.310 1513.990 2.680 ;
        RECT 1515.110 2.310 1530.550 2.680 ;
        RECT 1531.670 2.310 1547.110 2.680 ;
        RECT 1548.230 2.310 1563.670 2.680 ;
        RECT 1564.790 2.310 1580.230 2.680 ;
        RECT 1581.350 2.310 1596.790 2.680 ;
        RECT 1597.910 2.310 1613.350 2.680 ;
        RECT 1614.470 2.310 1629.910 2.680 ;
        RECT 1631.030 2.310 1647.390 2.680 ;
        RECT 1648.510 2.310 1663.950 2.680 ;
        RECT 1665.070 2.310 1680.510 2.680 ;
        RECT 1681.630 2.310 1697.070 2.680 ;
        RECT 1698.190 2.310 1713.630 2.680 ;
        RECT 1714.750 2.310 1730.190 2.680 ;
        RECT 1731.310 2.310 1746.750 2.680 ;
        RECT 1747.870 2.310 1763.310 2.680 ;
        RECT 1764.430 2.310 1779.870 2.680 ;
        RECT 1780.990 2.310 1796.430 2.680 ;
        RECT 1797.550 2.310 1812.990 2.680 ;
        RECT 1814.110 2.310 1830.470 2.680 ;
        RECT 1831.590 2.310 1847.030 2.680 ;
        RECT 1848.150 2.310 1863.590 2.680 ;
        RECT 1864.710 2.310 1880.150 2.680 ;
        RECT 1881.270 2.310 1896.710 2.680 ;
        RECT 1897.830 2.310 1913.270 2.680 ;
        RECT 1914.390 2.310 1929.830 2.680 ;
        RECT 1930.950 2.310 1946.390 2.680 ;
        RECT 1947.510 2.310 1962.950 2.680 ;
        RECT 1964.070 2.310 1979.510 2.680 ;
        RECT 1980.630 2.310 1996.070 2.680 ;
        RECT 1997.190 2.310 2013.550 2.680 ;
        RECT 2014.670 2.310 2030.110 2.680 ;
        RECT 2031.230 2.310 2046.670 2.680 ;
        RECT 2047.790 2.310 2063.230 2.680 ;
        RECT 2064.350 2.310 2079.790 2.680 ;
        RECT 2080.910 2.310 2096.350 2.680 ;
        RECT 2097.470 2.310 2112.910 2.680 ;
        RECT 2114.030 2.310 2129.470 2.680 ;
        RECT 2130.590 2.310 2146.030 2.680 ;
        RECT 2147.150 2.310 2162.590 2.680 ;
        RECT 2163.710 2.310 2179.150 2.680 ;
        RECT 2180.270 2.310 2196.630 2.680 ;
        RECT 2197.750 2.310 2213.190 2.680 ;
        RECT 2214.310 2.310 2229.750 2.680 ;
        RECT 2230.870 2.310 2246.310 2.680 ;
        RECT 2247.430 2.310 2262.870 2.680 ;
        RECT 2263.990 2.310 2279.430 2.680 ;
        RECT 2280.550 2.310 2295.990 2.680 ;
        RECT 2297.110 2.310 2312.550 2.680 ;
        RECT 2313.670 2.310 2329.110 2.680 ;
        RECT 2330.230 2.310 2345.670 2.680 ;
        RECT 2346.790 2.310 2362.230 2.680 ;
        RECT 2363.350 2.310 2379.710 2.680 ;
        RECT 2380.830 2.310 2396.270 2.680 ;
        RECT 2397.390 2.310 2412.830 2.680 ;
        RECT 2413.950 2.310 2429.390 2.680 ;
        RECT 2430.510 2.310 2445.950 2.680 ;
        RECT 2447.070 2.310 2462.510 2.680 ;
        RECT 2463.630 2.310 2479.070 2.680 ;
        RECT 2480.190 2.310 2495.630 2.680 ;
        RECT 2496.750 2.310 2512.190 2.680 ;
        RECT 2513.310 2.310 2528.750 2.680 ;
        RECT 2529.870 2.310 2545.310 2.680 ;
        RECT 2546.430 2.310 2562.790 2.680 ;
        RECT 2563.910 2.310 2579.350 2.680 ;
        RECT 2580.470 2.310 2595.910 2.680 ;
        RECT 2597.030 2.310 2612.470 2.680 ;
        RECT 2613.590 2.310 2629.030 2.680 ;
        RECT 2630.150 2.310 2645.590 2.680 ;
        RECT 2646.710 2.310 2662.150 2.680 ;
        RECT 2663.270 2.310 2678.710 2.680 ;
        RECT 2679.830 2.310 2695.270 2.680 ;
        RECT 2696.390 2.310 2711.830 2.680 ;
        RECT 2712.950 2.310 2728.390 2.680 ;
        RECT 2729.510 2.310 2745.870 2.680 ;
        RECT 2746.990 2.310 2762.430 2.680 ;
        RECT 2763.550 2.310 2778.990 2.680 ;
        RECT 2780.110 2.310 2795.550 2.680 ;
        RECT 2796.670 2.310 2812.110 2.680 ;
        RECT 2813.230 2.310 2828.670 2.680 ;
        RECT 2829.790 2.310 2845.230 2.680 ;
        RECT 2846.350 2.310 2861.790 2.680 ;
        RECT 2862.910 2.310 2878.350 2.680 ;
        RECT 2879.470 2.310 2894.910 2.680 ;
        RECT 2896.030 2.310 2911.470 2.680 ;
      LAYER met3 ;
        RECT 2.800 3517.660 2917.930 3518.825 ;
        RECT 2.400 3507.420 2917.930 3517.660 ;
        RECT 2.400 3505.420 2917.200 3507.420 ;
        RECT 2.400 3493.820 2917.930 3505.420 ;
        RECT 2.800 3491.820 2917.930 3493.820 ;
        RECT 2.400 3482.940 2917.930 3491.820 ;
        RECT 2.400 3480.940 2917.200 3482.940 ;
        RECT 2.400 3469.340 2917.930 3480.940 ;
        RECT 2.800 3467.340 2917.930 3469.340 ;
        RECT 2.400 3458.460 2917.930 3467.340 ;
        RECT 2.400 3456.460 2917.200 3458.460 ;
        RECT 2.400 3444.860 2917.930 3456.460 ;
        RECT 2.800 3442.860 2917.930 3444.860 ;
        RECT 2.400 3433.980 2917.930 3442.860 ;
        RECT 2.400 3431.980 2917.200 3433.980 ;
        RECT 2.400 3420.380 2917.930 3431.980 ;
        RECT 2.800 3418.380 2917.930 3420.380 ;
        RECT 2.400 3409.500 2917.930 3418.380 ;
        RECT 2.400 3407.500 2917.200 3409.500 ;
        RECT 2.400 3395.900 2917.930 3407.500 ;
        RECT 2.800 3393.900 2917.930 3395.900 ;
        RECT 2.400 3385.020 2917.930 3393.900 ;
        RECT 2.400 3383.020 2917.200 3385.020 ;
        RECT 2.400 3371.420 2917.930 3383.020 ;
        RECT 2.800 3369.420 2917.930 3371.420 ;
        RECT 2.400 3360.540 2917.930 3369.420 ;
        RECT 2.400 3358.540 2917.200 3360.540 ;
        RECT 2.400 3346.940 2917.930 3358.540 ;
        RECT 2.800 3344.940 2917.930 3346.940 ;
        RECT 2.400 3336.060 2917.930 3344.940 ;
        RECT 2.400 3334.060 2917.200 3336.060 ;
        RECT 2.400 3322.460 2917.930 3334.060 ;
        RECT 2.800 3320.460 2917.930 3322.460 ;
        RECT 2.400 3311.580 2917.930 3320.460 ;
        RECT 2.400 3309.580 2917.200 3311.580 ;
        RECT 2.400 3297.980 2917.930 3309.580 ;
        RECT 2.800 3295.980 2917.930 3297.980 ;
        RECT 2.400 3287.100 2917.930 3295.980 ;
        RECT 2.400 3285.100 2917.200 3287.100 ;
        RECT 2.400 3273.500 2917.930 3285.100 ;
        RECT 2.800 3271.500 2917.930 3273.500 ;
        RECT 2.400 3262.620 2917.930 3271.500 ;
        RECT 2.400 3260.620 2917.200 3262.620 ;
        RECT 2.400 3249.020 2917.930 3260.620 ;
        RECT 2.800 3247.020 2917.930 3249.020 ;
        RECT 2.400 3236.780 2917.930 3247.020 ;
        RECT 2.400 3234.780 2917.200 3236.780 ;
        RECT 2.400 3223.180 2917.930 3234.780 ;
        RECT 2.800 3221.180 2917.930 3223.180 ;
        RECT 2.400 3212.300 2917.930 3221.180 ;
        RECT 2.400 3210.300 2917.200 3212.300 ;
        RECT 2.400 3198.700 2917.930 3210.300 ;
        RECT 2.800 3196.700 2917.930 3198.700 ;
        RECT 2.400 3187.820 2917.930 3196.700 ;
        RECT 2.400 3185.820 2917.200 3187.820 ;
        RECT 2.400 3174.220 2917.930 3185.820 ;
        RECT 2.800 3172.220 2917.930 3174.220 ;
        RECT 2.400 3163.340 2917.930 3172.220 ;
        RECT 2.400 3161.340 2917.200 3163.340 ;
        RECT 2.400 3149.740 2917.930 3161.340 ;
        RECT 2.800 3147.740 2917.930 3149.740 ;
        RECT 2.400 3138.860 2917.930 3147.740 ;
        RECT 2.400 3136.860 2917.200 3138.860 ;
        RECT 2.400 3125.260 2917.930 3136.860 ;
        RECT 2.800 3123.260 2917.930 3125.260 ;
        RECT 2.400 3114.380 2917.930 3123.260 ;
        RECT 2.400 3112.380 2917.200 3114.380 ;
        RECT 2.400 3100.780 2917.930 3112.380 ;
        RECT 2.800 3098.780 2917.930 3100.780 ;
        RECT 2.400 3089.900 2917.930 3098.780 ;
        RECT 2.400 3087.900 2917.200 3089.900 ;
        RECT 2.400 3076.300 2917.930 3087.900 ;
        RECT 2.800 3074.300 2917.930 3076.300 ;
        RECT 2.400 3065.420 2917.930 3074.300 ;
        RECT 2.400 3063.420 2917.200 3065.420 ;
        RECT 2.400 3051.820 2917.930 3063.420 ;
        RECT 2.800 3049.820 2917.930 3051.820 ;
        RECT 2.400 3040.940 2917.930 3049.820 ;
        RECT 2.400 3038.940 2917.200 3040.940 ;
        RECT 2.400 3027.340 2917.930 3038.940 ;
        RECT 2.800 3025.340 2917.930 3027.340 ;
        RECT 2.400 3016.460 2917.930 3025.340 ;
        RECT 2.400 3014.460 2917.200 3016.460 ;
        RECT 2.400 3002.860 2917.930 3014.460 ;
        RECT 2.800 3000.860 2917.930 3002.860 ;
        RECT 2.400 2991.980 2917.930 3000.860 ;
        RECT 2.400 2989.980 2917.200 2991.980 ;
        RECT 2.400 2978.380 2917.930 2989.980 ;
        RECT 2.800 2976.380 2917.930 2978.380 ;
        RECT 2.400 2966.140 2917.930 2976.380 ;
        RECT 2.400 2964.140 2917.200 2966.140 ;
        RECT 2.400 2952.540 2917.930 2964.140 ;
        RECT 2.800 2950.540 2917.930 2952.540 ;
        RECT 2.400 2941.660 2917.930 2950.540 ;
        RECT 2.400 2939.660 2917.200 2941.660 ;
        RECT 2.400 2928.060 2917.930 2939.660 ;
        RECT 2.800 2926.060 2917.930 2928.060 ;
        RECT 2.400 2917.180 2917.930 2926.060 ;
        RECT 2.400 2915.180 2917.200 2917.180 ;
        RECT 2.400 2903.580 2917.930 2915.180 ;
        RECT 2.800 2901.580 2917.930 2903.580 ;
        RECT 2.400 2892.700 2917.930 2901.580 ;
        RECT 2.400 2890.700 2917.200 2892.700 ;
        RECT 2.400 2879.100 2917.930 2890.700 ;
        RECT 2.800 2877.100 2917.930 2879.100 ;
        RECT 2.400 2868.220 2917.930 2877.100 ;
        RECT 2.400 2866.220 2917.200 2868.220 ;
        RECT 2.400 2854.620 2917.930 2866.220 ;
        RECT 2.800 2852.620 2917.930 2854.620 ;
        RECT 2.400 2843.740 2917.930 2852.620 ;
        RECT 2.400 2841.740 2917.200 2843.740 ;
        RECT 2.400 2830.140 2917.930 2841.740 ;
        RECT 2.800 2828.140 2917.930 2830.140 ;
        RECT 2.400 2819.260 2917.930 2828.140 ;
        RECT 2.400 2817.260 2917.200 2819.260 ;
        RECT 2.400 2805.660 2917.930 2817.260 ;
        RECT 2.800 2803.660 2917.930 2805.660 ;
        RECT 2.400 2794.780 2917.930 2803.660 ;
        RECT 2.400 2792.780 2917.200 2794.780 ;
        RECT 2.400 2781.180 2917.930 2792.780 ;
        RECT 2.800 2779.180 2917.930 2781.180 ;
        RECT 2.400 2770.300 2917.930 2779.180 ;
        RECT 2.400 2768.300 2917.200 2770.300 ;
        RECT 2.400 2756.700 2917.930 2768.300 ;
        RECT 2.800 2754.700 2917.930 2756.700 ;
        RECT 2.400 2745.820 2917.930 2754.700 ;
        RECT 2.400 2743.820 2917.200 2745.820 ;
        RECT 2.400 2732.220 2917.930 2743.820 ;
        RECT 2.800 2730.220 2917.930 2732.220 ;
        RECT 2.400 2721.340 2917.930 2730.220 ;
        RECT 2.400 2719.340 2917.200 2721.340 ;
        RECT 2.400 2707.740 2917.930 2719.340 ;
        RECT 2.800 2705.740 2917.930 2707.740 ;
        RECT 2.400 2695.500 2917.930 2705.740 ;
        RECT 2.400 2693.500 2917.200 2695.500 ;
        RECT 2.400 2681.900 2917.930 2693.500 ;
        RECT 2.800 2679.900 2917.930 2681.900 ;
        RECT 2.400 2671.020 2917.930 2679.900 ;
        RECT 2.400 2669.020 2917.200 2671.020 ;
        RECT 2.400 2657.420 2917.930 2669.020 ;
        RECT 2.800 2655.420 2917.930 2657.420 ;
        RECT 2.400 2646.540 2917.930 2655.420 ;
        RECT 2.400 2644.540 2917.200 2646.540 ;
        RECT 2.400 2632.940 2917.930 2644.540 ;
        RECT 2.800 2630.940 2917.930 2632.940 ;
        RECT 2.400 2622.060 2917.930 2630.940 ;
        RECT 2.400 2620.060 2917.200 2622.060 ;
        RECT 2.400 2608.460 2917.930 2620.060 ;
        RECT 2.800 2606.460 2917.930 2608.460 ;
        RECT 2.400 2597.580 2917.930 2606.460 ;
        RECT 2.400 2595.580 2917.200 2597.580 ;
        RECT 2.400 2583.980 2917.930 2595.580 ;
        RECT 2.800 2581.980 2917.930 2583.980 ;
        RECT 2.400 2573.100 2917.930 2581.980 ;
        RECT 2.400 2571.100 2917.200 2573.100 ;
        RECT 2.400 2559.500 2917.930 2571.100 ;
        RECT 2.800 2557.500 2917.930 2559.500 ;
        RECT 2.400 2548.620 2917.930 2557.500 ;
        RECT 2.400 2546.620 2917.200 2548.620 ;
        RECT 2.400 2535.020 2917.930 2546.620 ;
        RECT 2.800 2533.020 2917.930 2535.020 ;
        RECT 2.400 2524.140 2917.930 2533.020 ;
        RECT 2.400 2522.140 2917.200 2524.140 ;
        RECT 2.400 2510.540 2917.930 2522.140 ;
        RECT 2.800 2508.540 2917.930 2510.540 ;
        RECT 2.400 2499.660 2917.930 2508.540 ;
        RECT 2.400 2497.660 2917.200 2499.660 ;
        RECT 2.400 2486.060 2917.930 2497.660 ;
        RECT 2.800 2484.060 2917.930 2486.060 ;
        RECT 2.400 2475.180 2917.930 2484.060 ;
        RECT 2.400 2473.180 2917.200 2475.180 ;
        RECT 2.400 2461.580 2917.930 2473.180 ;
        RECT 2.800 2459.580 2917.930 2461.580 ;
        RECT 2.400 2450.700 2917.930 2459.580 ;
        RECT 2.400 2448.700 2917.200 2450.700 ;
        RECT 2.400 2437.100 2917.930 2448.700 ;
        RECT 2.800 2435.100 2917.930 2437.100 ;
        RECT 2.400 2424.860 2917.930 2435.100 ;
        RECT 2.400 2422.860 2917.200 2424.860 ;
        RECT 2.400 2411.260 2917.930 2422.860 ;
        RECT 2.800 2409.260 2917.930 2411.260 ;
        RECT 2.400 2400.380 2917.930 2409.260 ;
        RECT 2.400 2398.380 2917.200 2400.380 ;
        RECT 2.400 2386.780 2917.930 2398.380 ;
        RECT 2.800 2384.780 2917.930 2386.780 ;
        RECT 2.400 2375.900 2917.930 2384.780 ;
        RECT 2.400 2373.900 2917.200 2375.900 ;
        RECT 2.400 2362.300 2917.930 2373.900 ;
        RECT 2.800 2360.300 2917.930 2362.300 ;
        RECT 2.400 2351.420 2917.930 2360.300 ;
        RECT 2.400 2349.420 2917.200 2351.420 ;
        RECT 2.400 2337.820 2917.930 2349.420 ;
        RECT 2.800 2335.820 2917.930 2337.820 ;
        RECT 2.400 2326.940 2917.930 2335.820 ;
        RECT 2.400 2324.940 2917.200 2326.940 ;
        RECT 2.400 2313.340 2917.930 2324.940 ;
        RECT 2.800 2311.340 2917.930 2313.340 ;
        RECT 2.400 2302.460 2917.930 2311.340 ;
        RECT 2.400 2300.460 2917.200 2302.460 ;
        RECT 2.400 2288.860 2917.930 2300.460 ;
        RECT 2.800 2286.860 2917.930 2288.860 ;
        RECT 2.400 2277.980 2917.930 2286.860 ;
        RECT 2.400 2275.980 2917.200 2277.980 ;
        RECT 2.400 2264.380 2917.930 2275.980 ;
        RECT 2.800 2262.380 2917.930 2264.380 ;
        RECT 2.400 2253.500 2917.930 2262.380 ;
        RECT 2.400 2251.500 2917.200 2253.500 ;
        RECT 2.400 2239.900 2917.930 2251.500 ;
        RECT 2.800 2237.900 2917.930 2239.900 ;
        RECT 2.400 2229.020 2917.930 2237.900 ;
        RECT 2.400 2227.020 2917.200 2229.020 ;
        RECT 2.400 2215.420 2917.930 2227.020 ;
        RECT 2.800 2213.420 2917.930 2215.420 ;
        RECT 2.400 2204.540 2917.930 2213.420 ;
        RECT 2.400 2202.540 2917.200 2204.540 ;
        RECT 2.400 2190.940 2917.930 2202.540 ;
        RECT 2.800 2188.940 2917.930 2190.940 ;
        RECT 2.400 2180.060 2917.930 2188.940 ;
        RECT 2.400 2178.060 2917.200 2180.060 ;
        RECT 2.400 2166.460 2917.930 2178.060 ;
        RECT 2.800 2164.460 2917.930 2166.460 ;
        RECT 2.400 2154.220 2917.930 2164.460 ;
        RECT 2.400 2152.220 2917.200 2154.220 ;
        RECT 2.400 2140.620 2917.930 2152.220 ;
        RECT 2.800 2138.620 2917.930 2140.620 ;
        RECT 2.400 2129.740 2917.930 2138.620 ;
        RECT 2.400 2127.740 2917.200 2129.740 ;
        RECT 2.400 2116.140 2917.930 2127.740 ;
        RECT 2.800 2114.140 2917.930 2116.140 ;
        RECT 2.400 2105.260 2917.930 2114.140 ;
        RECT 2.400 2103.260 2917.200 2105.260 ;
        RECT 2.400 2091.660 2917.930 2103.260 ;
        RECT 2.800 2089.660 2917.930 2091.660 ;
        RECT 2.400 2080.780 2917.930 2089.660 ;
        RECT 2.400 2078.780 2917.200 2080.780 ;
        RECT 2.400 2067.180 2917.930 2078.780 ;
        RECT 2.800 2065.180 2917.930 2067.180 ;
        RECT 2.400 2056.300 2917.930 2065.180 ;
        RECT 2.400 2054.300 2917.200 2056.300 ;
        RECT 2.400 2042.700 2917.930 2054.300 ;
        RECT 2.800 2040.700 2917.930 2042.700 ;
        RECT 2.400 2031.820 2917.930 2040.700 ;
        RECT 2.400 2029.820 2917.200 2031.820 ;
        RECT 2.400 2018.220 2917.930 2029.820 ;
        RECT 2.800 2016.220 2917.930 2018.220 ;
        RECT 2.400 2007.340 2917.930 2016.220 ;
        RECT 2.400 2005.340 2917.200 2007.340 ;
        RECT 2.400 1993.740 2917.930 2005.340 ;
        RECT 2.800 1991.740 2917.930 1993.740 ;
        RECT 2.400 1982.860 2917.930 1991.740 ;
        RECT 2.400 1980.860 2917.200 1982.860 ;
        RECT 2.400 1969.260 2917.930 1980.860 ;
        RECT 2.800 1967.260 2917.930 1969.260 ;
        RECT 2.400 1958.380 2917.930 1967.260 ;
        RECT 2.400 1956.380 2917.200 1958.380 ;
        RECT 2.400 1944.780 2917.930 1956.380 ;
        RECT 2.800 1942.780 2917.930 1944.780 ;
        RECT 2.400 1933.900 2917.930 1942.780 ;
        RECT 2.400 1931.900 2917.200 1933.900 ;
        RECT 2.400 1920.300 2917.930 1931.900 ;
        RECT 2.800 1918.300 2917.930 1920.300 ;
        RECT 2.400 1909.420 2917.930 1918.300 ;
        RECT 2.400 1907.420 2917.200 1909.420 ;
        RECT 2.400 1895.820 2917.930 1907.420 ;
        RECT 2.800 1893.820 2917.930 1895.820 ;
        RECT 2.400 1883.580 2917.930 1893.820 ;
        RECT 2.400 1881.580 2917.200 1883.580 ;
        RECT 2.400 1869.980 2917.930 1881.580 ;
        RECT 2.800 1867.980 2917.930 1869.980 ;
        RECT 2.400 1859.100 2917.930 1867.980 ;
        RECT 2.400 1857.100 2917.200 1859.100 ;
        RECT 2.400 1845.500 2917.930 1857.100 ;
        RECT 2.800 1843.500 2917.930 1845.500 ;
        RECT 2.400 1834.620 2917.930 1843.500 ;
        RECT 2.400 1832.620 2917.200 1834.620 ;
        RECT 2.400 1821.020 2917.930 1832.620 ;
        RECT 2.800 1819.020 2917.930 1821.020 ;
        RECT 2.400 1810.140 2917.930 1819.020 ;
        RECT 2.400 1808.140 2917.200 1810.140 ;
        RECT 2.400 1796.540 2917.930 1808.140 ;
        RECT 2.800 1794.540 2917.930 1796.540 ;
        RECT 2.400 1785.660 2917.930 1794.540 ;
        RECT 2.400 1783.660 2917.200 1785.660 ;
        RECT 2.400 1772.060 2917.930 1783.660 ;
        RECT 2.800 1770.060 2917.930 1772.060 ;
        RECT 2.400 1761.180 2917.930 1770.060 ;
        RECT 2.400 1759.180 2917.200 1761.180 ;
        RECT 2.400 1747.580 2917.930 1759.180 ;
        RECT 2.800 1745.580 2917.930 1747.580 ;
        RECT 2.400 1736.700 2917.930 1745.580 ;
        RECT 2.400 1734.700 2917.200 1736.700 ;
        RECT 2.400 1723.100 2917.930 1734.700 ;
        RECT 2.800 1721.100 2917.930 1723.100 ;
        RECT 2.400 1712.220 2917.930 1721.100 ;
        RECT 2.400 1710.220 2917.200 1712.220 ;
        RECT 2.400 1698.620 2917.930 1710.220 ;
        RECT 2.800 1696.620 2917.930 1698.620 ;
        RECT 2.400 1687.740 2917.930 1696.620 ;
        RECT 2.400 1685.740 2917.200 1687.740 ;
        RECT 2.400 1674.140 2917.930 1685.740 ;
        RECT 2.800 1672.140 2917.930 1674.140 ;
        RECT 2.400 1663.260 2917.930 1672.140 ;
        RECT 2.400 1661.260 2917.200 1663.260 ;
        RECT 2.400 1649.660 2917.930 1661.260 ;
        RECT 2.800 1647.660 2917.930 1649.660 ;
        RECT 2.400 1638.780 2917.930 1647.660 ;
        RECT 2.400 1636.780 2917.200 1638.780 ;
        RECT 2.400 1625.180 2917.930 1636.780 ;
        RECT 2.800 1623.180 2917.930 1625.180 ;
        RECT 2.400 1612.940 2917.930 1623.180 ;
        RECT 2.400 1610.940 2917.200 1612.940 ;
        RECT 2.400 1599.340 2917.930 1610.940 ;
        RECT 2.800 1597.340 2917.930 1599.340 ;
        RECT 2.400 1588.460 2917.930 1597.340 ;
        RECT 2.400 1586.460 2917.200 1588.460 ;
        RECT 2.400 1574.860 2917.930 1586.460 ;
        RECT 2.800 1572.860 2917.930 1574.860 ;
        RECT 2.400 1563.980 2917.930 1572.860 ;
        RECT 2.400 1561.980 2917.200 1563.980 ;
        RECT 2.400 1550.380 2917.930 1561.980 ;
        RECT 2.800 1548.380 2917.930 1550.380 ;
        RECT 2.400 1539.500 2917.930 1548.380 ;
        RECT 2.400 1537.500 2917.200 1539.500 ;
        RECT 2.400 1525.900 2917.930 1537.500 ;
        RECT 2.800 1523.900 2917.930 1525.900 ;
        RECT 2.400 1515.020 2917.930 1523.900 ;
        RECT 2.400 1513.020 2917.200 1515.020 ;
        RECT 2.400 1501.420 2917.930 1513.020 ;
        RECT 2.800 1499.420 2917.930 1501.420 ;
        RECT 2.400 1490.540 2917.930 1499.420 ;
        RECT 2.400 1488.540 2917.200 1490.540 ;
        RECT 2.400 1476.940 2917.930 1488.540 ;
        RECT 2.800 1474.940 2917.930 1476.940 ;
        RECT 2.400 1466.060 2917.930 1474.940 ;
        RECT 2.400 1464.060 2917.200 1466.060 ;
        RECT 2.400 1452.460 2917.930 1464.060 ;
        RECT 2.800 1450.460 2917.930 1452.460 ;
        RECT 2.400 1441.580 2917.930 1450.460 ;
        RECT 2.400 1439.580 2917.200 1441.580 ;
        RECT 2.400 1427.980 2917.930 1439.580 ;
        RECT 2.800 1425.980 2917.930 1427.980 ;
        RECT 2.400 1417.100 2917.930 1425.980 ;
        RECT 2.400 1415.100 2917.200 1417.100 ;
        RECT 2.400 1403.500 2917.930 1415.100 ;
        RECT 2.800 1401.500 2917.930 1403.500 ;
        RECT 2.400 1392.620 2917.930 1401.500 ;
        RECT 2.400 1390.620 2917.200 1392.620 ;
        RECT 2.400 1379.020 2917.930 1390.620 ;
        RECT 2.800 1377.020 2917.930 1379.020 ;
        RECT 2.400 1368.140 2917.930 1377.020 ;
        RECT 2.400 1366.140 2917.200 1368.140 ;
        RECT 2.400 1354.540 2917.930 1366.140 ;
        RECT 2.800 1352.540 2917.930 1354.540 ;
        RECT 2.400 1342.300 2917.930 1352.540 ;
        RECT 2.400 1340.300 2917.200 1342.300 ;
        RECT 2.400 1328.700 2917.930 1340.300 ;
        RECT 2.800 1326.700 2917.930 1328.700 ;
        RECT 2.400 1317.820 2917.930 1326.700 ;
        RECT 2.400 1315.820 2917.200 1317.820 ;
        RECT 2.400 1304.220 2917.930 1315.820 ;
        RECT 2.800 1302.220 2917.930 1304.220 ;
        RECT 2.400 1293.340 2917.930 1302.220 ;
        RECT 2.400 1291.340 2917.200 1293.340 ;
        RECT 2.400 1279.740 2917.930 1291.340 ;
        RECT 2.800 1277.740 2917.930 1279.740 ;
        RECT 2.400 1268.860 2917.930 1277.740 ;
        RECT 2.400 1266.860 2917.200 1268.860 ;
        RECT 2.400 1255.260 2917.930 1266.860 ;
        RECT 2.800 1253.260 2917.930 1255.260 ;
        RECT 2.400 1244.380 2917.930 1253.260 ;
        RECT 2.400 1242.380 2917.200 1244.380 ;
        RECT 2.400 1230.780 2917.930 1242.380 ;
        RECT 2.800 1228.780 2917.930 1230.780 ;
        RECT 2.400 1219.900 2917.930 1228.780 ;
        RECT 2.400 1217.900 2917.200 1219.900 ;
        RECT 2.400 1206.300 2917.930 1217.900 ;
        RECT 2.800 1204.300 2917.930 1206.300 ;
        RECT 2.400 1195.420 2917.930 1204.300 ;
        RECT 2.400 1193.420 2917.200 1195.420 ;
        RECT 2.400 1181.820 2917.930 1193.420 ;
        RECT 2.800 1179.820 2917.930 1181.820 ;
        RECT 2.400 1170.940 2917.930 1179.820 ;
        RECT 2.400 1168.940 2917.200 1170.940 ;
        RECT 2.400 1157.340 2917.930 1168.940 ;
        RECT 2.800 1155.340 2917.930 1157.340 ;
        RECT 2.400 1146.460 2917.930 1155.340 ;
        RECT 2.400 1144.460 2917.200 1146.460 ;
        RECT 2.400 1132.860 2917.930 1144.460 ;
        RECT 2.800 1130.860 2917.930 1132.860 ;
        RECT 2.400 1121.980 2917.930 1130.860 ;
        RECT 2.400 1119.980 2917.200 1121.980 ;
        RECT 2.400 1108.380 2917.930 1119.980 ;
        RECT 2.800 1106.380 2917.930 1108.380 ;
        RECT 2.400 1097.500 2917.930 1106.380 ;
        RECT 2.400 1095.500 2917.200 1097.500 ;
        RECT 2.400 1083.900 2917.930 1095.500 ;
        RECT 2.800 1081.900 2917.930 1083.900 ;
        RECT 2.400 1071.660 2917.930 1081.900 ;
        RECT 2.400 1069.660 2917.200 1071.660 ;
        RECT 2.400 1058.060 2917.930 1069.660 ;
        RECT 2.800 1056.060 2917.930 1058.060 ;
        RECT 2.400 1047.180 2917.930 1056.060 ;
        RECT 2.400 1045.180 2917.200 1047.180 ;
        RECT 2.400 1033.580 2917.930 1045.180 ;
        RECT 2.800 1031.580 2917.930 1033.580 ;
        RECT 2.400 1022.700 2917.930 1031.580 ;
        RECT 2.400 1020.700 2917.200 1022.700 ;
        RECT 2.400 1009.100 2917.930 1020.700 ;
        RECT 2.800 1007.100 2917.930 1009.100 ;
        RECT 2.400 998.220 2917.930 1007.100 ;
        RECT 2.400 996.220 2917.200 998.220 ;
        RECT 2.400 984.620 2917.930 996.220 ;
        RECT 2.800 982.620 2917.930 984.620 ;
        RECT 2.400 973.740 2917.930 982.620 ;
        RECT 2.400 971.740 2917.200 973.740 ;
        RECT 2.400 960.140 2917.930 971.740 ;
        RECT 2.800 958.140 2917.930 960.140 ;
        RECT 2.400 949.260 2917.930 958.140 ;
        RECT 2.400 947.260 2917.200 949.260 ;
        RECT 2.400 935.660 2917.930 947.260 ;
        RECT 2.800 933.660 2917.930 935.660 ;
        RECT 2.400 924.780 2917.930 933.660 ;
        RECT 2.400 922.780 2917.200 924.780 ;
        RECT 2.400 911.180 2917.930 922.780 ;
        RECT 2.800 909.180 2917.930 911.180 ;
        RECT 2.400 900.300 2917.930 909.180 ;
        RECT 2.400 898.300 2917.200 900.300 ;
        RECT 2.400 886.700 2917.930 898.300 ;
        RECT 2.800 884.700 2917.930 886.700 ;
        RECT 2.400 875.820 2917.930 884.700 ;
        RECT 2.400 873.820 2917.200 875.820 ;
        RECT 2.400 862.220 2917.930 873.820 ;
        RECT 2.800 860.220 2917.930 862.220 ;
        RECT 2.400 851.340 2917.930 860.220 ;
        RECT 2.400 849.340 2917.200 851.340 ;
        RECT 2.400 837.740 2917.930 849.340 ;
        RECT 2.800 835.740 2917.930 837.740 ;
        RECT 2.400 826.860 2917.930 835.740 ;
        RECT 2.400 824.860 2917.200 826.860 ;
        RECT 2.400 813.260 2917.930 824.860 ;
        RECT 2.800 811.260 2917.930 813.260 ;
        RECT 2.400 801.020 2917.930 811.260 ;
        RECT 2.400 799.020 2917.200 801.020 ;
        RECT 2.400 787.420 2917.930 799.020 ;
        RECT 2.800 785.420 2917.930 787.420 ;
        RECT 2.400 776.540 2917.930 785.420 ;
        RECT 2.400 774.540 2917.200 776.540 ;
        RECT 2.400 762.940 2917.930 774.540 ;
        RECT 2.800 760.940 2917.930 762.940 ;
        RECT 2.400 752.060 2917.930 760.940 ;
        RECT 2.400 750.060 2917.200 752.060 ;
        RECT 2.400 738.460 2917.930 750.060 ;
        RECT 2.800 736.460 2917.930 738.460 ;
        RECT 2.400 727.580 2917.930 736.460 ;
        RECT 2.400 725.580 2917.200 727.580 ;
        RECT 2.400 713.980 2917.930 725.580 ;
        RECT 2.800 711.980 2917.930 713.980 ;
        RECT 2.400 703.100 2917.930 711.980 ;
        RECT 2.400 701.100 2917.200 703.100 ;
        RECT 2.400 689.500 2917.930 701.100 ;
        RECT 2.800 687.500 2917.930 689.500 ;
        RECT 2.400 678.620 2917.930 687.500 ;
        RECT 2.400 676.620 2917.200 678.620 ;
        RECT 2.400 665.020 2917.930 676.620 ;
        RECT 2.800 663.020 2917.930 665.020 ;
        RECT 2.400 654.140 2917.930 663.020 ;
        RECT 2.400 652.140 2917.200 654.140 ;
        RECT 2.400 640.540 2917.930 652.140 ;
        RECT 2.800 638.540 2917.930 640.540 ;
        RECT 2.400 629.660 2917.930 638.540 ;
        RECT 2.400 627.660 2917.200 629.660 ;
        RECT 2.400 616.060 2917.930 627.660 ;
        RECT 2.800 614.060 2917.930 616.060 ;
        RECT 2.400 605.180 2917.930 614.060 ;
        RECT 2.400 603.180 2917.200 605.180 ;
        RECT 2.400 591.580 2917.930 603.180 ;
        RECT 2.800 589.580 2917.930 591.580 ;
        RECT 2.400 580.700 2917.930 589.580 ;
        RECT 2.400 578.700 2917.200 580.700 ;
        RECT 2.400 567.100 2917.930 578.700 ;
        RECT 2.800 565.100 2917.930 567.100 ;
        RECT 2.400 556.220 2917.930 565.100 ;
        RECT 2.400 554.220 2917.200 556.220 ;
        RECT 2.400 542.620 2917.930 554.220 ;
        RECT 2.800 540.620 2917.930 542.620 ;
        RECT 2.400 530.380 2917.930 540.620 ;
        RECT 2.400 528.380 2917.200 530.380 ;
        RECT 2.400 516.780 2917.930 528.380 ;
        RECT 2.800 514.780 2917.930 516.780 ;
        RECT 2.400 505.900 2917.930 514.780 ;
        RECT 2.400 503.900 2917.200 505.900 ;
        RECT 2.400 492.300 2917.930 503.900 ;
        RECT 2.800 490.300 2917.930 492.300 ;
        RECT 2.400 481.420 2917.930 490.300 ;
        RECT 2.400 479.420 2917.200 481.420 ;
        RECT 2.400 467.820 2917.930 479.420 ;
        RECT 2.800 465.820 2917.930 467.820 ;
        RECT 2.400 456.940 2917.930 465.820 ;
        RECT 2.400 454.940 2917.200 456.940 ;
        RECT 2.400 443.340 2917.930 454.940 ;
        RECT 2.800 441.340 2917.930 443.340 ;
        RECT 2.400 432.460 2917.930 441.340 ;
        RECT 2.400 430.460 2917.200 432.460 ;
        RECT 2.400 418.860 2917.930 430.460 ;
        RECT 2.800 416.860 2917.930 418.860 ;
        RECT 2.400 407.980 2917.930 416.860 ;
        RECT 2.400 405.980 2917.200 407.980 ;
        RECT 2.400 394.380 2917.930 405.980 ;
        RECT 2.800 392.380 2917.930 394.380 ;
        RECT 2.400 383.500 2917.930 392.380 ;
        RECT 2.400 381.500 2917.200 383.500 ;
        RECT 2.400 369.900 2917.930 381.500 ;
        RECT 2.800 367.900 2917.930 369.900 ;
        RECT 2.400 359.020 2917.930 367.900 ;
        RECT 2.400 357.020 2917.200 359.020 ;
        RECT 2.400 345.420 2917.930 357.020 ;
        RECT 2.800 343.420 2917.930 345.420 ;
        RECT 2.400 334.540 2917.930 343.420 ;
        RECT 2.400 332.540 2917.200 334.540 ;
        RECT 2.400 320.940 2917.930 332.540 ;
        RECT 2.800 318.940 2917.930 320.940 ;
        RECT 2.400 310.060 2917.930 318.940 ;
        RECT 2.400 308.060 2917.200 310.060 ;
        RECT 2.400 296.460 2917.930 308.060 ;
        RECT 2.800 294.460 2917.930 296.460 ;
        RECT 2.400 285.580 2917.930 294.460 ;
        RECT 2.400 283.580 2917.200 285.580 ;
        RECT 2.400 271.980 2917.930 283.580 ;
        RECT 2.800 269.980 2917.930 271.980 ;
        RECT 2.400 259.740 2917.930 269.980 ;
        RECT 2.400 257.740 2917.200 259.740 ;
        RECT 2.400 246.140 2917.930 257.740 ;
        RECT 2.800 244.140 2917.930 246.140 ;
        RECT 2.400 235.260 2917.930 244.140 ;
        RECT 2.400 233.260 2917.200 235.260 ;
        RECT 2.400 221.660 2917.930 233.260 ;
        RECT 2.800 219.660 2917.930 221.660 ;
        RECT 2.400 210.780 2917.930 219.660 ;
        RECT 2.400 208.780 2917.200 210.780 ;
        RECT 2.400 197.180 2917.930 208.780 ;
        RECT 2.800 195.180 2917.930 197.180 ;
        RECT 2.400 186.300 2917.930 195.180 ;
        RECT 2.400 184.300 2917.200 186.300 ;
        RECT 2.400 172.700 2917.930 184.300 ;
        RECT 2.800 170.700 2917.930 172.700 ;
        RECT 2.400 161.820 2917.930 170.700 ;
        RECT 2.400 159.820 2917.200 161.820 ;
        RECT 2.400 148.220 2917.930 159.820 ;
        RECT 2.800 146.220 2917.930 148.220 ;
        RECT 2.400 137.340 2917.930 146.220 ;
        RECT 2.400 135.340 2917.200 137.340 ;
        RECT 2.400 123.740 2917.930 135.340 ;
        RECT 2.800 121.740 2917.930 123.740 ;
        RECT 2.400 112.860 2917.930 121.740 ;
        RECT 2.400 110.860 2917.200 112.860 ;
        RECT 2.400 99.260 2917.930 110.860 ;
        RECT 2.800 97.260 2917.930 99.260 ;
        RECT 2.400 88.380 2917.930 97.260 ;
        RECT 2.400 86.380 2917.200 88.380 ;
        RECT 2.400 74.780 2917.930 86.380 ;
        RECT 2.800 72.780 2917.930 74.780 ;
        RECT 2.400 63.900 2917.930 72.780 ;
        RECT 2.400 61.900 2917.200 63.900 ;
        RECT 2.400 50.300 2917.930 61.900 ;
        RECT 2.800 48.300 2917.930 50.300 ;
        RECT 2.400 39.420 2917.930 48.300 ;
        RECT 2.400 37.420 2917.200 39.420 ;
        RECT 2.400 25.820 2917.930 37.420 ;
        RECT 2.800 23.820 2917.930 25.820 ;
        RECT 2.400 14.940 2917.930 23.820 ;
        RECT 2.400 13.775 2917.200 14.940 ;
      LAYER met4 ;
        RECT 194.415 14.455 2728.425 3505.225 ;
  END
END user_project_wrapper
END LIBRARY

