magic
tech sky130A
magscale 1 2
timestamp 1633664140
<< locali >>
rect 222301 663799 222335 664037
rect 382841 663799 382875 663901
rect 382691 663765 382875 663799
rect 41613 661351 41647 662337
rect 41463 661045 41889 661079
rect 39313 657271 39347 660773
rect 41429 660705 41521 660739
rect 40325 657067 40359 660501
rect 41429 657271 41463 660705
rect 42625 660263 42659 661249
rect 42717 660535 42751 662405
rect 49893 661079 49927 662609
rect 46121 660535 46155 660841
rect 46213 660739 46247 660841
rect 50939 660773 51181 660807
rect 46397 660671 46431 660773
rect 53021 660739 53055 660909
rect 59921 660875 59955 662609
rect 77217 661079 77251 662677
rect 110429 660943 110463 662677
rect 122481 661011 122515 663425
rect 153853 662235 153887 662337
rect 155233 661555 155267 662201
rect 155877 661555 155911 662065
rect 354045 660943 354079 662337
rect 358277 660875 358311 662337
rect 425069 661623 425103 662337
rect 427679 661521 427921 661555
rect 433901 661487 433935 662813
rect 479349 661147 479383 662813
rect 506397 661623 506431 662541
rect 515229 661011 515263 661657
rect 520197 661487 520231 661657
rect 541115 661181 541265 661215
rect 46305 660467 46339 660637
rect 46213 660263 46247 660433
rect 541909 654143 541943 660841
rect 543381 659515 543415 660229
rect 544117 659175 544151 660093
rect 544577 654823 544611 655605
rect 38945 650743 38979 652749
rect 542185 651287 542219 654313
rect 41429 45611 41463 50813
rect 40601 44387 40635 45577
rect 41797 43027 41831 45781
rect 541909 45557 541943 53805
rect 544669 45815 544703 46937
rect 540989 45523 541943 45557
rect 41981 44387 42015 44625
rect 41889 44183 41923 44353
rect 540989 44319 541023 45523
rect 541081 43163 541115 44285
rect 542277 43979 542311 44149
rect 541817 43639 541851 43809
rect 541725 43163 541759 43605
rect 542829 43571 542863 44625
rect 191849 42007 191883 42449
rect 436017 42007 436051 42449
rect 509157 42007 509191 42517
rect 536757 42007 536791 42585
rect 131129 38743 131163 40001
rect 542921 38879 542955 39457
rect 543013 39219 543047 39457
rect 536849 3451 536883 4029
rect 44281 3315 44315 3417
rect 44373 2839 44407 3281
rect 46949 3281 47133 3315
rect 46949 3247 46983 3281
rect 187743 3145 187893 3179
rect 59001 3077 59219 3111
rect 59001 3043 59035 3077
rect 59093 2907 59127 3009
rect 59185 2907 59219 3077
<< viali >>
rect 222301 664037 222335 664071
rect 382841 663901 382875 663935
rect 222301 663765 222335 663799
rect 382657 663765 382691 663799
rect 122481 663425 122515 663459
rect 77217 662677 77251 662711
rect 49893 662609 49927 662643
rect 42717 662405 42751 662439
rect 41613 662337 41647 662371
rect 41613 661317 41647 661351
rect 42625 661249 42659 661283
rect 41429 661045 41463 661079
rect 41889 661045 41923 661079
rect 39313 660773 39347 660807
rect 41521 660705 41555 660739
rect 39313 657237 39347 657271
rect 40325 660501 40359 660535
rect 49893 661045 49927 661079
rect 59921 662609 59955 662643
rect 53021 660909 53055 660943
rect 42717 660501 42751 660535
rect 46121 660841 46155 660875
rect 46213 660841 46247 660875
rect 46213 660705 46247 660739
rect 46397 660773 46431 660807
rect 50905 660773 50939 660807
rect 51181 660773 51215 660807
rect 77217 661045 77251 661079
rect 110429 662677 110463 662711
rect 433901 662813 433935 662847
rect 153853 662337 153887 662371
rect 354045 662337 354079 662371
rect 153853 662201 153887 662235
rect 155233 662201 155267 662235
rect 155233 661521 155267 661555
rect 155877 662065 155911 662099
rect 155877 661521 155911 661555
rect 122481 660977 122515 661011
rect 110429 660909 110463 660943
rect 354045 660909 354079 660943
rect 358277 662337 358311 662371
rect 59921 660841 59955 660875
rect 425069 662337 425103 662371
rect 425069 661589 425103 661623
rect 427645 661521 427679 661555
rect 427921 661521 427955 661555
rect 433901 661453 433935 661487
rect 479349 662813 479383 662847
rect 506397 662541 506431 662575
rect 506397 661589 506431 661623
rect 515229 661657 515263 661691
rect 479349 661113 479383 661147
rect 520197 661657 520231 661691
rect 520197 661453 520231 661487
rect 541081 661181 541115 661215
rect 541265 661181 541299 661215
rect 515229 660977 515263 661011
rect 358277 660841 358311 660875
rect 541909 660841 541943 660875
rect 53021 660705 53055 660739
rect 46121 660501 46155 660535
rect 46305 660637 46339 660671
rect 46397 660637 46431 660671
rect 42625 660229 42659 660263
rect 46213 660433 46247 660467
rect 46305 660433 46339 660467
rect 46213 660229 46247 660263
rect 41429 657237 41463 657271
rect 40325 657033 40359 657067
rect 543381 660229 543415 660263
rect 543381 659481 543415 659515
rect 544117 660093 544151 660127
rect 544117 659141 544151 659175
rect 544577 655605 544611 655639
rect 544577 654789 544611 654823
rect 541909 654109 541943 654143
rect 542185 654313 542219 654347
rect 38945 652749 38979 652783
rect 542185 651253 542219 651287
rect 38945 650709 38979 650743
rect 541909 53805 541943 53839
rect 41429 50813 41463 50847
rect 40601 45577 40635 45611
rect 41429 45577 41463 45611
rect 41797 45781 41831 45815
rect 40601 44353 40635 44387
rect 544669 46937 544703 46971
rect 544669 45781 544703 45815
rect 41981 44625 42015 44659
rect 41889 44353 41923 44387
rect 41981 44353 42015 44387
rect 542829 44625 542863 44659
rect 540989 44285 541023 44319
rect 541081 44285 541115 44319
rect 41889 44149 41923 44183
rect 542277 44149 542311 44183
rect 542277 43945 542311 43979
rect 541817 43809 541851 43843
rect 541081 43129 541115 43163
rect 541725 43605 541759 43639
rect 541817 43605 541851 43639
rect 542829 43537 542863 43571
rect 541725 43129 541759 43163
rect 41797 42993 41831 43027
rect 536757 42585 536791 42619
rect 509157 42517 509191 42551
rect 191849 42449 191883 42483
rect 191849 41973 191883 42007
rect 436017 42449 436051 42483
rect 436017 41973 436051 42007
rect 509157 41973 509191 42007
rect 536757 41973 536791 42007
rect 131129 40001 131163 40035
rect 542921 39457 542955 39491
rect 543013 39457 543047 39491
rect 543013 39185 543047 39219
rect 542921 38845 542955 38879
rect 131129 38709 131163 38743
rect 536849 4029 536883 4063
rect 44281 3417 44315 3451
rect 536849 3417 536883 3451
rect 44281 3281 44315 3315
rect 44373 3281 44407 3315
rect 47133 3281 47167 3315
rect 46949 3213 46983 3247
rect 187709 3145 187743 3179
rect 187893 3145 187927 3179
rect 59001 3009 59035 3043
rect 59093 3009 59127 3043
rect 59093 2873 59127 2907
rect 59185 2873 59219 2907
rect 44373 2805 44407 2839
<< metal1 >>
rect 314654 702992 314660 703044
rect 314712 703032 314718 703044
rect 315942 703032 315948 703044
rect 314712 703004 315948 703032
rect 314712 702992 314718 703004
rect 315942 702992 315948 703004
rect 316000 702992 316006 703044
rect 3418 702448 3424 702500
rect 3476 702488 3482 702500
rect 7742 702488 7748 702500
rect 3476 702460 7748 702488
rect 3476 702448 3482 702460
rect 7742 702448 7748 702460
rect 7800 702448 7806 702500
rect 38654 700952 38660 701004
rect 38712 700992 38718 701004
rect 73062 700992 73068 701004
rect 38712 700964 73068 700992
rect 38712 700952 38718 700964
rect 73062 700952 73068 700964
rect 73120 700952 73126 701004
rect 73154 700952 73160 701004
rect 73212 700992 73218 701004
rect 575566 700992 575572 701004
rect 73212 700964 575572 700992
rect 73212 700952 73218 700964
rect 575566 700952 575572 700964
rect 575624 700952 575630 701004
rect 40034 700884 40040 700936
rect 40092 700924 40098 700936
rect 239398 700924 239404 700936
rect 40092 700896 239404 700924
rect 40092 700884 40098 700896
rect 239398 700884 239404 700896
rect 239456 700884 239462 700936
rect 302694 700884 302700 700936
rect 302752 700924 302758 700936
rect 543918 700924 543924 700936
rect 302752 700896 543924 700924
rect 302752 700884 302758 700896
rect 543918 700884 543924 700896
rect 543976 700884 543982 700936
rect 38010 700816 38016 700868
rect 38068 700856 38074 700868
rect 276014 700856 276020 700868
rect 38068 700828 276020 700856
rect 38068 700816 38074 700828
rect 276014 700816 276020 700828
rect 276072 700816 276078 700868
rect 299382 700816 299388 700868
rect 299440 700856 299446 700868
rect 541986 700856 541992 700868
rect 299440 700828 541992 700856
rect 299440 700816 299446 700828
rect 541986 700816 541992 700828
rect 542044 700816 542050 700868
rect 37090 700748 37096 700800
rect 37148 700788 37154 700800
rect 312630 700788 312636 700800
rect 37148 700760 312636 700788
rect 37148 700748 37154 700760
rect 312630 700748 312636 700760
rect 312688 700748 312694 700800
rect 329374 700748 329380 700800
rect 329432 700788 329438 700800
rect 543826 700788 543832 700800
rect 329432 700760 543832 700788
rect 329432 700748 329438 700760
rect 543826 700748 543832 700760
rect 543884 700748 543890 700800
rect 41874 700680 41880 700732
rect 41932 700720 41938 700732
rect 56318 700720 56324 700732
rect 41932 700692 56324 700720
rect 41932 700680 41938 700692
rect 56318 700680 56324 700692
rect 56376 700680 56382 700732
rect 62942 700680 62948 700732
rect 63000 700720 63006 700732
rect 352466 700720 352472 700732
rect 63000 700692 352472 700720
rect 63000 700680 63006 700692
rect 352466 700680 352472 700692
rect 352524 700680 352530 700732
rect 352742 700680 352748 700732
rect 352800 700720 352806 700732
rect 385862 700720 385868 700732
rect 352800 700692 385868 700720
rect 352800 700680 352806 700692
rect 385862 700680 385868 700692
rect 385920 700680 385926 700732
rect 398742 700680 398748 700732
rect 398800 700720 398806 700732
rect 415854 700720 415860 700732
rect 398800 700692 415860 700720
rect 398800 700680 398806 700692
rect 415854 700680 415860 700692
rect 415912 700680 415918 700732
rect 419166 700680 419172 700732
rect 419224 700720 419230 700732
rect 542262 700720 542268 700732
rect 419224 700692 542268 700720
rect 419224 700680 419230 700692
rect 542262 700680 542268 700692
rect 542320 700680 542326 700732
rect 38102 700612 38108 700664
rect 38160 700652 38166 700664
rect 335998 700652 336004 700664
rect 38160 700624 336004 700652
rect 38160 700612 38166 700624
rect 335998 700612 336004 700624
rect 336056 700612 336062 700664
rect 345934 700612 345940 700664
rect 345992 700652 345998 700664
rect 543734 700652 543740 700664
rect 345992 700624 543740 700652
rect 345992 700612 345998 700624
rect 543734 700612 543740 700624
rect 543792 700612 543798 700664
rect 38838 700544 38844 700596
rect 38896 700584 38902 700596
rect 362494 700584 362500 700596
rect 38896 700556 362500 700584
rect 38896 700544 38902 700556
rect 362494 700544 362500 700556
rect 362552 700544 362558 700596
rect 395798 700544 395804 700596
rect 395856 700584 395862 700596
rect 543642 700584 543648 700596
rect 395856 700556 543648 700584
rect 395856 700544 395862 700556
rect 543642 700544 543648 700556
rect 543700 700544 543706 700596
rect 37458 700476 37464 700528
rect 37516 700516 37522 700528
rect 149606 700516 149612 700528
rect 37516 700488 149612 700516
rect 37516 700476 37522 700488
rect 149606 700476 149612 700488
rect 149664 700476 149670 700528
rect 166166 700476 166172 700528
rect 166224 700516 166230 700528
rect 542814 700516 542820 700528
rect 166224 700488 542820 700516
rect 166224 700476 166230 700488
rect 542814 700476 542820 700488
rect 542872 700476 542878 700528
rect 39942 700408 39948 700460
rect 40000 700448 40006 700460
rect 422478 700448 422484 700460
rect 40000 700420 422484 700448
rect 40000 700408 40006 700420
rect 422478 700408 422484 700420
rect 422536 700408 422542 700460
rect 455782 700408 455788 700460
rect 455840 700448 455846 700460
rect 542170 700448 542176 700460
rect 455840 700420 542176 700448
rect 455840 700408 455846 700420
rect 542170 700408 542176 700420
rect 542228 700408 542234 700460
rect 547414 700408 547420 700460
rect 547472 700448 547478 700460
rect 555694 700448 555700 700460
rect 547472 700420 555700 700448
rect 547472 700408 547478 700420
rect 555694 700408 555700 700420
rect 555752 700408 555758 700460
rect 39666 700340 39672 700392
rect 39724 700380 39730 700392
rect 432414 700380 432420 700392
rect 39724 700352 432420 700380
rect 39724 700340 39730 700352
rect 432414 700340 432420 700352
rect 432472 700340 432478 700392
rect 459462 700340 459468 700392
rect 459520 700380 459526 700392
rect 578878 700380 578884 700392
rect 459520 700352 578884 700380
rect 459520 700340 459526 700352
rect 578878 700340 578884 700352
rect 578936 700340 578942 700392
rect 38286 700272 38292 700324
rect 38344 700312 38350 700324
rect 495710 700312 495716 700324
rect 38344 700284 495716 700312
rect 38344 700272 38350 700284
rect 495710 700272 495716 700284
rect 495768 700272 495774 700324
rect 508958 700272 508964 700324
rect 509016 700312 509022 700324
rect 544194 700312 544200 700324
rect 509016 700284 544200 700312
rect 509016 700272 509022 700284
rect 544194 700272 544200 700284
rect 544252 700272 544258 700324
rect 550174 700272 550180 700324
rect 550232 700312 550238 700324
rect 562318 700312 562324 700324
rect 550232 700284 562324 700312
rect 550232 700272 550238 700284
rect 562318 700272 562324 700284
rect 562376 700272 562382 700324
rect 39482 700204 39488 700256
rect 39540 700244 39546 700256
rect 216030 700244 216036 700256
rect 39540 700216 216036 700244
rect 39540 700204 39546 700216
rect 216030 700204 216036 700216
rect 216088 700204 216094 700256
rect 236086 700204 236092 700256
rect 236144 700244 236150 700256
rect 242158 700244 242164 700256
rect 236144 700216 242164 700244
rect 236144 700204 236150 700216
rect 242158 700204 242164 700216
rect 242216 700204 242222 700256
rect 282638 700204 282644 700256
rect 282696 700244 282702 700256
rect 491938 700244 491944 700256
rect 282696 700216 491944 700244
rect 282696 700204 282702 700216
rect 491938 700204 491944 700216
rect 491996 700204 492002 700256
rect 40402 700136 40408 700188
rect 40460 700176 40466 700188
rect 189534 700176 189540 700188
rect 40460 700148 189540 700176
rect 40460 700136 40466 700148
rect 189534 700136 189540 700148
rect 189592 700136 189598 700188
rect 256142 700136 256148 700188
rect 256200 700176 256206 700188
rect 324314 700176 324320 700188
rect 256200 700148 324320 700176
rect 256200 700136 256206 700148
rect 324314 700136 324320 700148
rect 324372 700136 324378 700188
rect 325602 700136 325608 700188
rect 325660 700176 325666 700188
rect 462406 700176 462412 700188
rect 325660 700148 462412 700176
rect 325660 700136 325666 700148
rect 462406 700136 462412 700148
rect 462464 700136 462470 700188
rect 464982 700136 464988 700188
rect 465040 700176 465046 700188
rect 535638 700176 535644 700188
rect 465040 700148 535644 700176
rect 465040 700136 465046 700148
rect 535638 700136 535644 700148
rect 535696 700136 535702 700188
rect 9766 700068 9772 700120
rect 9824 700108 9830 700120
rect 10962 700108 10968 700120
rect 9824 700080 10968 700108
rect 9824 700068 9830 700080
rect 10962 700068 10968 700080
rect 11020 700068 11026 700120
rect 26326 700068 26332 700120
rect 26384 700108 26390 700120
rect 27522 700108 27528 700120
rect 26384 700080 27528 700108
rect 26384 700068 26390 700080
rect 27522 700068 27528 700080
rect 27580 700068 27586 700120
rect 41598 700068 41604 700120
rect 41656 700108 41662 700120
rect 146294 700108 146300 700120
rect 41656 700080 146300 700108
rect 41656 700068 41662 700080
rect 146294 700068 146300 700080
rect 146352 700068 146358 700120
rect 169478 700068 169484 700120
rect 169536 700108 169542 700120
rect 175918 700108 175924 700120
rect 169536 700080 175924 700108
rect 169536 700068 169542 700080
rect 175918 700068 175924 700080
rect 175976 700068 175982 700120
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 326798 700108 326804 700120
rect 202840 700080 326804 700108
rect 202840 700068 202846 700080
rect 326798 700068 326804 700080
rect 326856 700068 326862 700120
rect 352650 700068 352656 700120
rect 352708 700108 352714 700120
rect 382550 700108 382556 700120
rect 352708 700080 382556 700108
rect 352708 700068 352714 700080
rect 382550 700068 382556 700080
rect 382608 700068 382614 700120
rect 416038 700068 416044 700120
rect 416096 700108 416102 700120
rect 429102 700108 429108 700120
rect 416096 700080 429108 700108
rect 416096 700068 416102 700080
rect 429102 700068 429108 700080
rect 429160 700068 429166 700120
rect 461578 700068 461584 700120
rect 461636 700108 461642 700120
rect 479150 700108 479156 700120
rect 461636 700080 479156 700108
rect 461636 700068 461642 700080
rect 479150 700068 479156 700080
rect 479208 700068 479214 700120
rect 485774 700068 485780 700120
rect 485832 700108 485838 700120
rect 542906 700108 542912 700120
rect 485832 700080 542912 700108
rect 485832 700068 485838 700080
rect 542906 700068 542912 700080
rect 542964 700068 542970 700120
rect 41230 700000 41236 700052
rect 41288 700040 41294 700052
rect 139486 700040 139492 700052
rect 41288 700012 139492 700040
rect 41288 700000 41294 700012
rect 139486 700000 139492 700012
rect 139544 700000 139550 700052
rect 152918 700000 152924 700052
rect 152976 700040 152982 700052
rect 264974 700040 264980 700052
rect 152976 700012 264980 700040
rect 152976 700000 152982 700012
rect 264974 700000 264980 700012
rect 265032 700000 265038 700052
rect 489178 700000 489184 700052
rect 489236 700040 489242 700052
rect 499022 700040 499028 700052
rect 489236 700012 499028 700040
rect 489236 700000 489242 700012
rect 499022 700000 499028 700012
rect 499080 700000 499086 700052
rect 39206 699932 39212 699984
rect 39264 699972 39270 699984
rect 39264 699944 45554 699972
rect 39264 699932 39270 699944
rect 38378 699864 38384 699916
rect 38436 699904 38442 699916
rect 43070 699904 43076 699916
rect 38436 699876 43076 699904
rect 38436 699864 38442 699876
rect 43070 699864 43076 699876
rect 43128 699864 43134 699916
rect 45526 699904 45554 699944
rect 54478 699932 54484 699984
rect 54536 699972 54542 699984
rect 159542 699972 159548 699984
rect 54536 699944 159548 699972
rect 54536 699932 54542 699944
rect 159542 699932 159548 699944
rect 159600 699932 159606 699984
rect 425790 699932 425796 699984
rect 425848 699972 425854 699984
rect 426342 699972 426348 699984
rect 425848 699944 426348 699972
rect 425848 699932 425854 699944
rect 426342 699932 426348 699944
rect 426400 699932 426406 699984
rect 132862 699904 132868 699916
rect 45526 699876 132868 699904
rect 132862 699864 132868 699876
rect 132920 699864 132926 699916
rect 150342 699864 150348 699916
rect 150400 699904 150406 699916
rect 206094 699904 206100 699916
rect 150400 699876 206100 699904
rect 150400 699864 150406 699876
rect 206094 699864 206100 699876
rect 206152 699864 206158 699916
rect 36446 699796 36452 699848
rect 36504 699836 36510 699848
rect 37182 699836 37188 699848
rect 36504 699808 37188 699836
rect 36504 699796 36510 699808
rect 37182 699796 37188 699808
rect 37240 699796 37246 699848
rect 41046 699796 41052 699848
rect 41104 699836 41110 699848
rect 106182 699836 106188 699848
rect 41104 699808 106188 699836
rect 41104 699796 41110 699808
rect 106182 699796 106188 699808
rect 106240 699796 106246 699848
rect 112990 699796 112996 699848
rect 113048 699836 113054 699848
rect 128998 699836 129004 699848
rect 113048 699808 129004 699836
rect 113048 699796 113054 699808
rect 128998 699796 129004 699808
rect 129056 699796 129062 699848
rect 142798 699796 142804 699848
rect 142856 699836 142862 699848
rect 152458 699836 152464 699848
rect 142856 699808 152464 699836
rect 142856 699796 142862 699808
rect 152458 699796 152464 699808
rect 152516 699796 152522 699848
rect 3142 699728 3148 699780
rect 3200 699768 3206 699780
rect 6178 699768 6184 699780
rect 3200 699740 6184 699768
rect 3200 699728 3206 699740
rect 6178 699728 6184 699740
rect 6236 699728 6242 699780
rect 41322 699728 41328 699780
rect 41380 699768 41386 699780
rect 41380 699740 76328 699768
rect 41380 699728 41386 699740
rect 19702 699660 19708 699712
rect 19760 699700 19766 699712
rect 20622 699700 20628 699712
rect 19760 699672 20628 699700
rect 19760 699660 19766 699672
rect 20622 699660 20628 699672
rect 20680 699660 20686 699712
rect 41782 699660 41788 699712
rect 41840 699700 41846 699712
rect 46382 699700 46388 699712
rect 41840 699672 46388 699700
rect 41840 699660 41846 699672
rect 46382 699660 46388 699672
rect 46440 699660 46446 699712
rect 53006 699660 53012 699712
rect 53064 699700 53070 699712
rect 53650 699700 53656 699712
rect 53064 699672 53656 699700
rect 53064 699660 53070 699672
rect 53650 699660 53656 699672
rect 53708 699660 53714 699712
rect 66898 699660 66904 699712
rect 66956 699700 66962 699712
rect 66956 699672 69520 699700
rect 66956 699660 66962 699672
rect 69492 699632 69520 699672
rect 69566 699660 69572 699712
rect 69624 699700 69630 699712
rect 70302 699700 70308 699712
rect 69624 699672 70308 699700
rect 69624 699660 69630 699672
rect 70302 699660 70308 699672
rect 70360 699660 70366 699712
rect 70412 699672 76236 699700
rect 70412 699632 70440 699672
rect 69492 699604 70440 699632
rect 76208 699564 76236 699672
rect 76300 699632 76328 699740
rect 76374 699728 76380 699780
rect 76432 699768 76438 699780
rect 77202 699768 77208 699780
rect 76432 699740 77208 699768
rect 76432 699728 76438 699740
rect 77202 699728 77208 699740
rect 77260 699728 77266 699780
rect 82998 699768 83004 699780
rect 77312 699740 83004 699768
rect 77312 699632 77340 699740
rect 82998 699728 83004 699740
rect 83056 699728 83062 699780
rect 86310 699728 86316 699780
rect 86368 699768 86374 699780
rect 86862 699768 86868 699780
rect 86368 699740 86868 699768
rect 86368 699728 86374 699740
rect 86862 699728 86868 699740
rect 86920 699728 86926 699780
rect 102870 699728 102876 699780
rect 102928 699768 102934 699780
rect 109678 699768 109684 699780
rect 102928 699740 109684 699768
rect 102928 699728 102934 699740
rect 109678 699728 109684 699740
rect 109736 699728 109742 699780
rect 180058 699728 180064 699780
rect 180116 699768 180122 699780
rect 182910 699768 182916 699780
rect 180116 699740 182916 699768
rect 180116 699728 180122 699740
rect 182910 699728 182916 699740
rect 182968 699728 182974 699780
rect 99558 699700 99564 699712
rect 76300 699604 77340 699632
rect 77404 699672 99564 699700
rect 77404 699564 77432 699672
rect 99558 699660 99564 699672
rect 99616 699660 99622 699712
rect 119614 699660 119620 699712
rect 119672 699700 119678 699712
rect 122098 699700 122104 699712
rect 119672 699672 122104 699700
rect 119672 699660 119678 699672
rect 122098 699660 122104 699672
rect 122156 699660 122162 699712
rect 122926 699660 122932 699712
rect 122984 699700 122990 699712
rect 124122 699700 124128 699712
rect 122984 699672 124128 699700
rect 122984 699660 122990 699672
rect 124122 699660 124128 699672
rect 124180 699660 124186 699712
rect 172790 699660 172796 699712
rect 172848 699700 172854 699712
rect 173802 699700 173808 699712
rect 172848 699672 173808 699700
rect 172848 699660 172854 699672
rect 173802 699660 173808 699672
rect 173860 699660 173866 699712
rect 179414 699660 179420 699712
rect 179472 699700 179478 699712
rect 180702 699700 180708 699712
rect 179472 699672 180708 699700
rect 179472 699660 179478 699672
rect 180702 699660 180708 699672
rect 180760 699660 180766 699712
rect 196158 699660 196164 699712
rect 196216 699700 196222 699712
rect 197262 699700 197268 699712
rect 196216 699672 197268 699700
rect 196216 699660 196222 699672
rect 197262 699660 197268 699672
rect 197320 699660 197326 699712
rect 199470 699660 199476 699712
rect 199528 699700 199534 699712
rect 200022 699700 200028 699712
rect 199528 699672 200028 699700
rect 199528 699660 199534 699672
rect 200022 699660 200028 699672
rect 200080 699660 200086 699712
rect 212718 699660 212724 699712
rect 212776 699700 212782 699712
rect 213822 699700 213828 699712
rect 212776 699672 213828 699700
rect 212776 699660 212782 699672
rect 213822 699660 213828 699672
rect 213880 699660 213886 699712
rect 219526 699660 219532 699712
rect 219584 699700 219590 699712
rect 220722 699700 220728 699712
rect 219584 699672 220728 699700
rect 219584 699660 219590 699672
rect 220722 699660 220728 699672
rect 220780 699660 220786 699712
rect 222838 699660 222844 699712
rect 222896 699700 222902 699712
rect 223482 699700 223488 699712
rect 222896 699672 223488 699700
rect 222896 699660 222902 699672
rect 223482 699660 223488 699672
rect 223540 699660 223546 699712
rect 259454 699660 259460 699712
rect 259512 699700 259518 699712
rect 260742 699700 260748 699712
rect 259512 699672 260748 699700
rect 259512 699660 259518 699672
rect 260742 699660 260748 699672
rect 260800 699660 260806 699712
rect 269390 699660 269396 699712
rect 269448 699700 269454 699712
rect 270402 699700 270408 699712
rect 269448 699672 270408 699700
rect 269448 699660 269454 699672
rect 270402 699660 270408 699672
rect 270460 699660 270466 699712
rect 272702 699660 272708 699712
rect 272760 699700 272766 699712
rect 273162 699700 273168 699712
rect 272760 699672 273168 699700
rect 272760 699660 272766 699672
rect 273162 699660 273168 699672
rect 273220 699660 273226 699712
rect 278774 699660 278780 699712
rect 278832 699700 278838 699712
rect 279326 699700 279332 699712
rect 278832 699672 279332 699700
rect 278832 699660 278838 699672
rect 279326 699660 279332 699672
rect 279384 699660 279390 699712
rect 289262 699660 289268 699712
rect 289320 699700 289326 699712
rect 289722 699700 289728 699712
rect 289320 699672 289728 699700
rect 289320 699660 289326 699672
rect 289722 699660 289728 699672
rect 289780 699660 289786 699712
rect 309318 699660 309324 699712
rect 309376 699700 309382 699712
rect 310422 699700 310428 699712
rect 309376 699672 310428 699700
rect 309376 699660 309382 699672
rect 310422 699660 310428 699672
rect 310480 699660 310486 699712
rect 352558 699660 352564 699712
rect 352616 699700 352622 699712
rect 353202 699700 353208 699712
rect 352616 699672 353208 699700
rect 352616 699660 352622 699672
rect 353202 699660 353208 699672
rect 353260 699660 353266 699712
rect 436738 699660 436744 699712
rect 436796 699700 436802 699712
rect 439222 699700 439228 699712
rect 436796 699672 439228 699700
rect 436796 699660 436802 699672
rect 439222 699660 439228 699672
rect 439280 699660 439286 699712
rect 465718 699660 465724 699712
rect 465776 699700 465782 699712
rect 466362 699700 466368 699712
rect 465776 699672 466368 699700
rect 465776 699660 465782 699672
rect 466362 699660 466368 699672
rect 466420 699660 466426 699712
rect 505646 699660 505652 699712
rect 505704 699700 505710 699712
rect 506382 699700 506388 699712
rect 505704 699672 506388 699700
rect 505704 699660 505710 699672
rect 506382 699660 506388 699672
rect 506440 699660 506446 699712
rect 512638 699660 512644 699712
rect 512696 699700 512702 699712
rect 515766 699700 515772 699712
rect 512696 699672 515772 699700
rect 512696 699660 512702 699672
rect 515766 699660 515772 699672
rect 515824 699660 515830 699712
rect 519078 699660 519084 699712
rect 519136 699700 519142 699712
rect 520182 699700 520188 699712
rect 519136 699672 520188 699700
rect 519136 699660 519142 699672
rect 520182 699660 520188 699672
rect 520240 699660 520246 699712
rect 326798 699592 326804 699644
rect 326856 699632 326862 699644
rect 334618 699632 334624 699644
rect 326856 699604 334624 699632
rect 326856 699592 326862 699604
rect 334618 699592 334624 699604
rect 334676 699592 334682 699644
rect 76208 699536 77432 699564
rect 29638 698912 29644 698964
rect 29696 698952 29702 698964
rect 59998 698952 60004 698964
rect 29696 698924 60004 698952
rect 29696 698912 29702 698924
rect 59998 698912 60004 698924
rect 60056 698912 60062 698964
rect 68554 698912 68560 698964
rect 68612 698952 68618 698964
rect 129550 698952 129556 698964
rect 68612 698924 129556 698952
rect 68612 698912 68618 698924
rect 129550 698912 129556 698924
rect 129608 698912 129614 698964
rect 264974 698640 264980 698692
rect 265032 698680 265038 698692
rect 266998 698680 267004 698692
rect 265032 698652 267004 698680
rect 265032 698640 265038 698652
rect 266998 698640 267004 698652
rect 267056 698640 267062 698692
rect 3234 698300 3240 698352
rect 3292 698340 3298 698352
rect 509878 698340 509884 698352
rect 3292 698312 509884 698340
rect 3292 698300 3298 698312
rect 509878 698300 509884 698312
rect 509936 698300 509942 698352
rect 64138 697552 64144 697604
rect 64196 697592 64202 697604
rect 68554 697592 68560 697604
rect 64196 697564 68560 697592
rect 64196 697552 64202 697564
rect 68554 697552 68560 697564
rect 68612 697552 68618 697604
rect 244918 697552 244924 697604
rect 244976 697592 244982 697604
rect 262766 697592 262772 697604
rect 244976 697564 262772 697592
rect 244976 697552 244982 697564
rect 262766 697552 262772 697564
rect 262824 697552 262830 697604
rect 285950 697552 285956 697604
rect 286008 697592 286014 697604
rect 294598 697592 294604 697604
rect 286008 697564 294604 697592
rect 286008 697552 286014 697564
rect 294598 697552 294604 697564
rect 294656 697552 294662 697604
rect 109770 696192 109776 696244
rect 109828 696232 109834 696244
rect 135898 696232 135904 696244
rect 109828 696204 135904 696232
rect 109828 696192 109834 696204
rect 135898 696192 135904 696204
rect 135956 696192 135962 696244
rect 324314 696192 324320 696244
rect 324372 696232 324378 696244
rect 331858 696232 331864 696244
rect 324372 696204 331864 696232
rect 324372 696192 324378 696204
rect 331858 696192 331864 696204
rect 331916 696192 331922 696244
rect 3142 692792 3148 692844
rect 3200 692832 3206 692844
rect 10318 692832 10324 692844
rect 3200 692804 10324 692832
rect 3200 692792 3206 692804
rect 10318 692792 10324 692804
rect 10376 692792 10382 692844
rect 294598 692724 294604 692776
rect 294656 692764 294662 692776
rect 298002 692764 298008 692776
rect 294656 692736 298008 692764
rect 294656 692724 294662 692736
rect 298002 692724 298008 692736
rect 298060 692724 298066 692776
rect 334618 692588 334624 692640
rect 334676 692628 334682 692640
rect 336458 692628 336464 692640
rect 334676 692600 336464 692628
rect 334676 692588 334682 692600
rect 336458 692588 336464 692600
rect 336516 692588 336522 692640
rect 544838 691364 544844 691416
rect 544896 691404 544902 691416
rect 580166 691404 580172 691416
rect 544896 691376 580172 691404
rect 544896 691364 544902 691376
rect 580166 691364 580172 691376
rect 580224 691364 580230 691416
rect 331858 690004 331864 690056
rect 331916 690044 331922 690056
rect 333238 690044 333244 690056
rect 331916 690016 333244 690044
rect 331916 690004 331922 690016
rect 333238 690004 333244 690016
rect 333296 690004 333302 690056
rect 336458 689732 336464 689784
rect 336516 689772 336522 689784
rect 338758 689772 338764 689784
rect 336516 689744 338764 689772
rect 336516 689732 336522 689744
rect 338758 689732 338764 689744
rect 338816 689732 338822 689784
rect 298002 688984 298008 689036
rect 298060 689024 298066 689036
rect 305086 689024 305092 689036
rect 298060 688996 305092 689024
rect 298060 688984 298066 688996
rect 305086 688984 305092 688996
rect 305144 688984 305150 689036
rect 62758 687420 62764 687472
rect 62816 687460 62822 687472
rect 64138 687460 64144 687472
rect 62816 687432 64144 687460
rect 62816 687420 62822 687432
rect 64138 687420 64144 687432
rect 64196 687420 64202 687472
rect 266998 686468 267004 686520
rect 267056 686508 267062 686520
rect 273254 686508 273260 686520
rect 267056 686480 273260 686508
rect 267056 686468 267062 686480
rect 273254 686468 273260 686480
rect 273312 686468 273318 686520
rect 552750 685856 552756 685908
rect 552808 685896 552814 685908
rect 579614 685896 579620 685908
rect 552808 685868 579620 685896
rect 552808 685856 552814 685868
rect 579614 685856 579620 685868
rect 579672 685856 579678 685908
rect 234522 685108 234528 685160
rect 234580 685148 234586 685160
rect 244918 685148 244924 685160
rect 234580 685120 244924 685148
rect 234580 685108 234586 685120
rect 244918 685108 244924 685120
rect 244976 685108 244982 685160
rect 305086 685108 305092 685160
rect 305144 685148 305150 685160
rect 310238 685148 310244 685160
rect 305144 685120 310244 685148
rect 305144 685108 305150 685120
rect 310238 685108 310244 685120
rect 310296 685108 310302 685160
rect 273254 684496 273260 684548
rect 273312 684536 273318 684548
rect 273312 684508 277394 684536
rect 273312 684496 273318 684508
rect 277366 684468 277394 684508
rect 278866 684468 278872 684480
rect 277366 684440 278872 684468
rect 278866 684428 278872 684440
rect 278924 684428 278930 684480
rect 310238 682592 310244 682644
rect 310296 682632 310302 682644
rect 318702 682632 318708 682644
rect 310296 682604 318708 682632
rect 310296 682592 310302 682604
rect 318702 682592 318708 682604
rect 318760 682592 318766 682644
rect 278866 681708 278872 681760
rect 278924 681748 278930 681760
rect 280798 681748 280804 681760
rect 278924 681720 280804 681748
rect 278924 681708 278930 681720
rect 280798 681708 280804 681720
rect 280856 681708 280862 681760
rect 338758 681708 338764 681760
rect 338816 681748 338822 681760
rect 340138 681748 340144 681760
rect 338816 681720 340144 681748
rect 338816 681708 338822 681720
rect 340138 681708 340144 681720
rect 340196 681708 340202 681760
rect 333238 680892 333244 680944
rect 333296 680932 333302 680944
rect 333974 680932 333980 680944
rect 333296 680904 333980 680932
rect 333296 680892 333302 680904
rect 333974 680892 333980 680904
rect 334032 680892 334038 680944
rect 332502 680348 332508 680400
rect 332560 680388 332566 680400
rect 580166 680388 580172 680400
rect 332560 680360 580172 680388
rect 332560 680348 332566 680360
rect 580166 680348 580172 680360
rect 580224 680348 580230 680400
rect 318702 679600 318708 679652
rect 318760 679640 318766 679652
rect 331858 679640 331864 679652
rect 318760 679612 331864 679640
rect 318760 679600 318766 679612
rect 331858 679600 331864 679612
rect 331916 679600 331922 679652
rect 61286 678988 61292 679040
rect 61344 679028 61350 679040
rect 62758 679028 62764 679040
rect 61344 679000 62764 679028
rect 61344 678988 61350 679000
rect 62758 678988 62764 679000
rect 62816 678988 62822 679040
rect 228358 678240 228364 678292
rect 228416 678280 228422 678292
rect 234522 678280 234528 678292
rect 228416 678252 234528 678280
rect 228416 678240 228422 678252
rect 234522 678240 234528 678252
rect 234580 678240 234586 678292
rect 333974 676812 333980 676864
rect 334032 676852 334038 676864
rect 341518 676852 341524 676864
rect 334032 676824 341524 676852
rect 334032 676812 334038 676824
rect 341518 676812 341524 676824
rect 341576 676812 341582 676864
rect 171870 676336 171876 676388
rect 171928 676376 171934 676388
rect 175274 676376 175280 676388
rect 171928 676348 175280 676376
rect 171928 676336 171934 676348
rect 175274 676336 175280 676348
rect 175332 676336 175338 676388
rect 59722 675792 59728 675844
rect 59780 675832 59786 675844
rect 61286 675832 61292 675844
rect 59780 675804 61292 675832
rect 59780 675792 59786 675804
rect 61286 675792 61292 675804
rect 61344 675792 61350 675844
rect 166258 673480 166264 673532
rect 166316 673520 166322 673532
rect 171870 673520 171876 673532
rect 166316 673492 171876 673520
rect 166316 673480 166322 673492
rect 171870 673480 171876 673492
rect 171928 673480 171934 673532
rect 341518 672528 341524 672580
rect 341576 672568 341582 672580
rect 346302 672568 346308 672580
rect 341576 672540 346308 672568
rect 341576 672528 341582 672540
rect 346302 672528 346308 672540
rect 346360 672528 346366 672580
rect 280798 672052 280804 672104
rect 280856 672092 280862 672104
rect 280856 672064 281580 672092
rect 280856 672052 280862 672064
rect 281552 672024 281580 672064
rect 282914 672024 282920 672036
rect 281552 671996 282920 672024
rect 282914 671984 282920 671996
rect 282972 671984 282978 672036
rect 331858 671304 331864 671356
rect 331916 671344 331922 671356
rect 343634 671344 343640 671356
rect 331916 671316 343640 671344
rect 331916 671304 331922 671316
rect 343634 671304 343640 671316
rect 343692 671304 343698 671356
rect 554038 670692 554044 670744
rect 554096 670732 554102 670744
rect 580166 670732 580172 670744
rect 554096 670704 580172 670732
rect 554096 670692 554102 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 340138 669332 340144 669384
rect 340196 669372 340202 669384
rect 340196 669344 345014 669372
rect 340196 669332 340202 669344
rect 344986 669236 345014 669344
rect 346118 669236 346124 669248
rect 344986 669208 346124 669236
rect 346118 669196 346124 669208
rect 346176 669196 346182 669248
rect 282914 668584 282920 668636
rect 282972 668624 282978 668636
rect 284938 668624 284944 668636
rect 282972 668596 284944 668624
rect 282972 668584 282978 668596
rect 284938 668584 284944 668596
rect 284996 668584 285002 668636
rect 222102 668108 222108 668160
rect 222160 668148 222166 668160
rect 228358 668148 228364 668160
rect 222160 668120 228364 668148
rect 222160 668108 222166 668120
rect 228358 668108 228364 668120
rect 228416 668108 228422 668160
rect 57790 666544 57796 666596
rect 57848 666584 57854 666596
rect 59722 666584 59728 666596
rect 57848 666556 59728 666584
rect 57848 666544 57854 666556
rect 59722 666544 59728 666556
rect 59780 666544 59786 666596
rect 548518 666544 548524 666596
rect 548576 666584 548582 666596
rect 579614 666584 579620 666596
rect 548576 666556 579620 666584
rect 548576 666544 548582 666556
rect 579614 666544 579620 666556
rect 579672 666544 579678 666596
rect 64874 666476 64880 666528
rect 64932 666516 64938 666528
rect 66898 666516 66904 666528
rect 64932 666488 66904 666516
rect 64932 666476 64938 666488
rect 66898 666476 66904 666488
rect 66956 666476 66962 666528
rect 98178 666476 98184 666528
rect 98236 666516 98242 666528
rect 252554 666516 252560 666528
rect 98236 666488 252560 666516
rect 98236 666476 98242 666488
rect 252554 666476 252560 666488
rect 252612 666476 252618 666528
rect 270402 666476 270408 666528
rect 270460 666516 270466 666528
rect 388806 666516 388812 666528
rect 270460 666488 388812 666516
rect 270460 666476 270466 666488
rect 388806 666476 388812 666488
rect 388864 666476 388870 666528
rect 161842 666408 161848 666460
rect 161900 666448 161906 666460
rect 325694 666448 325700 666460
rect 161900 666420 325700 666448
rect 161900 666408 161906 666420
rect 325694 666408 325700 666420
rect 325752 666408 325758 666460
rect 340506 666408 340512 666460
rect 340564 666448 340570 666460
rect 352742 666448 352748 666460
rect 340564 666420 352748 666448
rect 340564 666408 340570 666420
rect 352742 666408 352748 666420
rect 352800 666408 352806 666460
rect 353202 666408 353208 666460
rect 353260 666448 353266 666460
rect 428182 666448 428188 666460
rect 353260 666420 428188 666448
rect 353260 666408 353266 666420
rect 428182 666408 428188 666420
rect 428240 666408 428246 666460
rect 197262 666340 197268 666392
rect 197320 666380 197326 666392
rect 407114 666380 407120 666392
rect 197320 666352 407120 666380
rect 197320 666340 197326 666352
rect 407114 666340 407120 666352
rect 407172 666340 407178 666392
rect 70946 666272 70952 666324
rect 71004 666312 71010 666324
rect 292574 666312 292580 666324
rect 71004 666284 292580 666312
rect 71004 666272 71010 666284
rect 292574 666272 292580 666284
rect 292632 666272 292638 666324
rect 316218 666272 316224 666324
rect 316276 666312 316282 666324
rect 441614 666312 441620 666324
rect 316276 666284 441620 666312
rect 316276 666272 316282 666284
rect 441614 666272 441620 666284
rect 441672 666272 441678 666324
rect 136542 666204 136548 666256
rect 136600 666244 136606 666256
rect 358630 666244 358636 666256
rect 136600 666216 358636 666244
rect 136600 666204 136606 666216
rect 358630 666204 358636 666216
rect 358688 666204 358694 666256
rect 422202 666204 422208 666256
rect 422260 666244 422266 666256
rect 436738 666244 436744 666256
rect 422260 666216 436744 666244
rect 422260 666204 422266 666216
rect 436738 666204 436744 666216
rect 436796 666204 436802 666256
rect 122098 666136 122104 666188
rect 122156 666176 122162 666188
rect 146478 666176 146484 666188
rect 122156 666148 146484 666176
rect 122156 666136 122162 666148
rect 146478 666136 146484 666148
rect 146536 666136 146542 666188
rect 164786 666136 164792 666188
rect 164844 666176 164850 666188
rect 481634 666176 481640 666188
rect 164844 666148 481640 666176
rect 164844 666136 164850 666148
rect 481634 666136 481640 666148
rect 481692 666136 481698 666188
rect 79962 666068 79968 666120
rect 80020 666108 80026 666120
rect 431310 666108 431316 666120
rect 80020 666080 431316 666108
rect 80020 666068 80026 666080
rect 431310 666068 431316 666080
rect 431368 666068 431374 666120
rect 492214 666068 492220 666120
rect 492272 666108 492278 666120
rect 512638 666108 512644 666120
rect 492272 666080 512644 666108
rect 492272 666068 492278 666080
rect 512638 666068 512644 666080
rect 512696 666068 512702 666120
rect 124122 666000 124128 666052
rect 124180 666040 124186 666052
rect 510062 666040 510068 666052
rect 124180 666012 510068 666040
rect 124180 666000 124186 666012
rect 510062 666000 510068 666012
rect 510120 666000 510126 666052
rect 86034 665932 86040 665984
rect 86092 665972 86098 665984
rect 95234 665972 95240 665984
rect 86092 665944 95240 665972
rect 86092 665932 86098 665944
rect 95234 665932 95240 665944
rect 95292 665932 95298 665984
rect 134426 665932 134432 665984
rect 134484 665972 134490 665984
rect 531314 665972 531320 665984
rect 134484 665944 531320 665972
rect 134484 665932 134490 665944
rect 531314 665932 531320 665944
rect 531372 665932 531378 665984
rect 39574 665864 39580 665916
rect 39632 665904 39638 665916
rect 519078 665904 519084 665916
rect 39632 665876 519084 665904
rect 39632 665864 39638 665876
rect 519078 665864 519084 665876
rect 519136 665864 519142 665916
rect 52730 665796 52736 665848
rect 52788 665836 52794 665848
rect 552014 665836 552020 665848
rect 52788 665808 552020 665836
rect 52788 665796 52794 665808
rect 552014 665796 552020 665808
rect 552072 665796 552078 665848
rect 167914 665728 167920 665780
rect 167972 665768 167978 665780
rect 318794 665768 318800 665780
rect 167972 665740 318800 665768
rect 167972 665728 167978 665740
rect 318794 665728 318800 665740
rect 318852 665728 318858 665780
rect 346394 665728 346400 665780
rect 346452 665768 346458 665780
rect 349062 665768 349068 665780
rect 346452 665740 349068 665768
rect 346452 665728 346458 665740
rect 349062 665728 349068 665740
rect 349120 665728 349126 665780
rect 86862 665660 86868 665712
rect 86920 665700 86926 665712
rect 207198 665700 207204 665712
rect 86920 665672 207204 665700
rect 86920 665660 86926 665672
rect 207198 665660 207204 665672
rect 207256 665660 207262 665712
rect 223482 665660 223488 665712
rect 223540 665700 223546 665712
rect 246574 665700 246580 665712
rect 223540 665672 246580 665700
rect 223540 665660 223546 665672
rect 246574 665660 246580 665672
rect 246632 665660 246638 665712
rect 193122 665592 193128 665644
rect 193180 665632 193186 665644
rect 231302 665632 231308 665644
rect 193180 665604 231308 665632
rect 193180 665592 193186 665604
rect 231302 665592 231308 665604
rect 231360 665592 231366 665644
rect 214650 665184 214656 665236
rect 214708 665224 214714 665236
rect 222102 665224 222108 665236
rect 214708 665196 222108 665224
rect 214708 665184 214714 665196
rect 222102 665184 222108 665196
rect 222160 665184 222166 665236
rect 49786 665116 49792 665168
rect 49844 665156 49850 665168
rect 54478 665156 54484 665168
rect 49844 665128 54484 665156
rect 49844 665116 49850 665128
rect 54478 665116 54484 665128
rect 54536 665116 54542 665168
rect 113266 665116 113272 665168
rect 113324 665156 113330 665168
rect 539594 665156 539600 665168
rect 113324 665128 539600 665156
rect 113324 665116 113330 665128
rect 539594 665116 539600 665128
rect 539652 665116 539658 665168
rect 5166 665048 5172 665100
rect 5224 665088 5230 665100
rect 101030 665088 101036 665100
rect 5224 665060 101036 665088
rect 5224 665048 5230 665060
rect 101030 665048 101036 665060
rect 101088 665048 101094 665100
rect 107194 665048 107200 665100
rect 107252 665088 107258 665100
rect 551278 665088 551284 665100
rect 107252 665060 551284 665088
rect 107252 665048 107258 665060
rect 551278 665048 551284 665060
rect 551336 665048 551342 665100
rect 38562 664980 38568 665032
rect 38620 665020 38626 665032
rect 46566 665020 46572 665032
rect 38620 664992 46572 665020
rect 38620 664980 38626 664992
rect 46566 664980 46572 664992
rect 46624 664980 46630 665032
rect 59998 664980 60004 665032
rect 60056 665020 60062 665032
rect 104158 665020 104164 665032
rect 60056 664992 104164 665020
rect 60056 664980 60062 664992
rect 104158 664980 104164 664992
rect 104216 664980 104222 665032
rect 135898 664980 135904 665032
rect 135956 665020 135962 665032
rect 140406 665020 140412 665032
rect 135956 664992 140412 665020
rect 135956 664980 135962 664992
rect 140406 664980 140412 664992
rect 140464 664980 140470 665032
rect 176930 664980 176936 665032
rect 176988 665020 176994 665032
rect 180058 665020 180064 665032
rect 176988 664992 180064 665020
rect 176988 664980 176994 664992
rect 180058 664980 180064 664992
rect 180116 664980 180122 665032
rect 249702 664980 249708 665032
rect 249760 665020 249766 665032
rect 252554 665020 252560 665032
rect 249760 664992 252560 665020
rect 249760 664980 249766 664992
rect 252554 664980 252560 664992
rect 252612 664980 252618 665032
rect 266262 664980 266268 665032
rect 266320 665020 266326 665032
rect 276750 665020 276756 665032
rect 266320 664992 276756 665020
rect 266320 664980 266326 664992
rect 276750 664980 276756 664992
rect 276808 664980 276814 665032
rect 304074 664980 304080 665032
rect 304132 665020 304138 665032
rect 304994 665020 305000 665032
rect 304132 664992 305000 665020
rect 304132 664980 304138 664992
rect 304994 664980 305000 664992
rect 305052 664980 305058 665032
rect 331306 664980 331312 665032
rect 331364 665020 331370 665032
rect 332502 665020 332508 665032
rect 331364 664992 332508 665020
rect 331364 664980 331370 664992
rect 332502 664980 332508 664992
rect 332560 664980 332566 665032
rect 337378 664980 337384 665032
rect 337436 665020 337442 665032
rect 342254 665020 342260 665032
rect 337436 664992 342260 665020
rect 337436 664980 337442 664992
rect 342254 664980 342260 664992
rect 342312 664980 342318 665032
rect 373810 664980 373816 665032
rect 373868 665020 373874 665032
rect 389174 665020 389180 665032
rect 373868 664992 389180 665020
rect 373868 664980 373874 664992
rect 389174 664980 389180 664992
rect 389232 664980 389238 665032
rect 413186 664980 413192 665032
rect 413244 665020 413250 665032
rect 416038 665020 416044 665032
rect 413244 664992 416044 665020
rect 413244 664980 413250 664992
rect 416038 664980 416044 664992
rect 416096 664980 416102 665032
rect 458634 664980 458640 665032
rect 458692 665020 458698 665032
rect 459462 665020 459468 665032
rect 458692 664992 459468 665020
rect 458692 664980 458698 664992
rect 459462 664980 459468 664992
rect 459520 664980 459526 665032
rect 473722 664980 473728 665032
rect 473780 665020 473786 665032
rect 489178 665020 489184 665032
rect 473780 664992 489184 665020
rect 473780 664980 473786 664992
rect 489178 664980 489184 664992
rect 489236 664980 489242 665032
rect 491938 664980 491944 665032
rect 491996 665020 492002 665032
rect 500954 665020 500960 665032
rect 491996 664992 500960 665020
rect 491996 664980 492002 664992
rect 500954 664980 500960 664992
rect 501012 664980 501018 665032
rect 509878 664980 509884 665032
rect 509936 665020 509942 665032
rect 516134 665020 516140 665032
rect 509936 664992 516140 665020
rect 509936 664980 509942 664992
rect 516134 664980 516140 664992
rect 516192 664980 516198 665032
rect 10594 664912 10600 664964
rect 10652 664952 10658 664964
rect 61654 664952 61660 664964
rect 10652 664924 61660 664952
rect 10652 664912 10658 664924
rect 61654 664912 61660 664924
rect 61712 664912 61718 664964
rect 70302 664912 70308 664964
rect 70360 664952 70366 664964
rect 219158 664952 219164 664964
rect 70360 664924 219164 664952
rect 70360 664912 70366 664924
rect 219158 664912 219164 664924
rect 219216 664912 219222 664964
rect 234522 664912 234528 664964
rect 234580 664952 234586 664964
rect 352650 664952 352656 664964
rect 234580 664924 352656 664952
rect 234580 664912 234586 664924
rect 352650 664912 352656 664924
rect 352708 664912 352714 664964
rect 361666 664912 361672 664964
rect 361724 664952 361730 664964
rect 368474 664952 368480 664964
rect 361724 664924 368480 664952
rect 361724 664912 361730 664924
rect 368474 664912 368480 664924
rect 368532 664912 368538 664964
rect 385954 664912 385960 664964
rect 386012 664952 386018 664964
rect 401594 664952 401600 664964
rect 386012 664924 401600 664952
rect 386012 664912 386018 664924
rect 401594 664912 401600 664924
rect 401652 664912 401658 664964
rect 466362 664912 466368 664964
rect 466420 664952 466426 664964
rect 531314 664952 531320 664964
rect 466420 664924 531320 664952
rect 466420 664912 466426 664924
rect 531314 664912 531320 664924
rect 531372 664912 531378 664964
rect 7926 664844 7932 664896
rect 7984 664884 7990 664896
rect 79870 664884 79876 664896
rect 7984 664856 79876 664884
rect 7984 664844 7990 664856
rect 79870 664844 79876 664856
rect 79928 664844 79934 664896
rect 89622 664844 89628 664896
rect 89680 664884 89686 664896
rect 270678 664884 270684 664896
rect 89680 664856 270684 664884
rect 89680 664844 89686 664856
rect 270678 664844 270684 664856
rect 270736 664844 270742 664896
rect 289722 664844 289728 664896
rect 289780 664884 289786 664896
rect 470686 664884 470692 664896
rect 289780 664856 470692 664884
rect 289780 664844 289786 664856
rect 470686 664844 470692 664856
rect 470744 664844 470750 664896
rect 482922 664844 482928 664896
rect 482980 664884 482986 664896
rect 553026 664884 553032 664896
rect 482980 664856 553032 664884
rect 482980 664844 482986 664856
rect 553026 664844 553032 664856
rect 553084 664844 553090 664896
rect 5074 664776 5080 664828
rect 5132 664816 5138 664828
rect 82998 664816 83004 664828
rect 5132 664788 83004 664816
rect 5132 664776 5138 664788
rect 82998 664776 83004 664788
rect 83056 664776 83062 664828
rect 119338 664776 119344 664828
rect 119396 664816 119402 664828
rect 314654 664816 314660 664828
rect 119396 664788 314660 664816
rect 119396 664776 119402 664788
rect 314654 664776 314660 664788
rect 314712 664776 314718 664828
rect 352558 664776 352564 664828
rect 352616 664816 352622 664828
rect 443454 664816 443460 664828
rect 352616 664788 443460 664816
rect 352616 664776 352622 664788
rect 443454 664776 443460 664788
rect 443512 664776 443518 664828
rect 446490 664776 446496 664828
rect 446548 664816 446554 664828
rect 542354 664816 542360 664828
rect 446548 664788 542360 664816
rect 446548 664776 446554 664788
rect 542354 664776 542360 664788
rect 542412 664776 542418 664828
rect 27522 664708 27528 664760
rect 27580 664748 27586 664760
rect 225230 664748 225236 664760
rect 27580 664720 225236 664748
rect 27580 664708 27586 664720
rect 225230 664708 225236 664720
rect 225288 664708 225294 664760
rect 242158 664708 242164 664760
rect 242216 664748 242222 664760
rect 258534 664748 258540 664760
rect 242216 664720 258540 664748
rect 242216 664708 242222 664720
rect 258534 664708 258540 664720
rect 258592 664708 258598 664760
rect 273162 664708 273168 664760
rect 273220 664748 273226 664760
rect 282914 664748 282920 664760
rect 273220 664720 282920 664748
rect 273220 664708 273226 664720
rect 282914 664708 282920 664720
rect 282972 664708 282978 664760
rect 334434 664708 334440 664760
rect 334492 664748 334498 664760
rect 521654 664748 521660 664760
rect 334492 664720 521660 664748
rect 334492 664708 334498 664720
rect 521654 664708 521660 664720
rect 521712 664708 521718 664760
rect 522298 664708 522304 664760
rect 522356 664748 522362 664760
rect 547598 664748 547604 664760
rect 522356 664720 547604 664748
rect 522356 664708 522362 664720
rect 547598 664708 547604 664720
rect 547656 664708 547662 664760
rect 9582 664640 9588 664692
rect 9640 664680 9646 664692
rect 89070 664680 89076 664692
rect 9640 664652 89076 664680
rect 9640 664640 9646 664652
rect 89070 664640 89076 664652
rect 89128 664640 89134 664692
rect 109678 664640 109684 664692
rect 109736 664680 109742 664692
rect 125318 664680 125324 664692
rect 109736 664652 125324 664680
rect 109736 664640 109742 664652
rect 125318 664640 125324 664652
rect 125376 664640 125382 664692
rect 128998 664640 129004 664692
rect 129056 664680 129062 664692
rect 137462 664680 137468 664692
rect 129056 664652 137468 664680
rect 129056 664640 129062 664652
rect 137462 664640 137468 664652
rect 137520 664640 137526 664692
rect 189074 664640 189080 664692
rect 189132 664680 189138 664692
rect 458174 664680 458180 664692
rect 189132 664652 458180 664680
rect 189132 664640 189138 664652
rect 458174 664640 458180 664652
rect 458232 664640 458238 664692
rect 476850 664640 476856 664692
rect 476908 664680 476914 664692
rect 548886 664680 548892 664692
rect 476908 664652 548892 664680
rect 476908 664640 476914 664652
rect 548886 664640 548892 664652
rect 548944 664640 548950 664692
rect 3418 664572 3424 664624
rect 3476 664612 3482 664624
rect 143534 664612 143540 664624
rect 3476 664584 143540 664612
rect 3476 664572 3482 664584
rect 143534 664572 143540 664584
rect 143592 664572 143598 664624
rect 152458 664572 152464 664624
rect 152516 664612 152522 664624
rect 170766 664612 170772 664624
rect 152516 664584 170772 664612
rect 152516 664572 152522 664584
rect 170766 664572 170772 664584
rect 170824 664572 170830 664624
rect 182910 664612 182916 664624
rect 175936 664584 182916 664612
rect 10870 664504 10876 664556
rect 10928 664544 10934 664556
rect 173710 664544 173716 664556
rect 10928 664516 173716 664544
rect 10928 664504 10934 664516
rect 173710 664504 173716 664516
rect 173768 664504 173774 664556
rect 9306 664436 9312 664488
rect 9364 664476 9370 664488
rect 175936 664476 175964 664584
rect 182910 664572 182916 664584
rect 182968 664572 182974 664624
rect 455506 664572 455512 664624
rect 455564 664612 455570 664624
rect 461578 664612 461584 664624
rect 455564 664584 461584 664612
rect 455564 664572 455570 664584
rect 461578 664572 461584 664584
rect 461636 664572 461642 664624
rect 485866 664572 485872 664624
rect 485924 664612 485930 664624
rect 551370 664612 551376 664624
rect 485924 664584 551376 664612
rect 485924 664572 485930 664584
rect 551370 664572 551376 664584
rect 551428 664572 551434 664624
rect 176010 664504 176016 664556
rect 176068 664544 176074 664556
rect 185854 664544 185860 664556
rect 176068 664516 185860 664544
rect 176068 664504 176074 664516
rect 185854 664504 185860 664516
rect 185912 664504 185918 664556
rect 186222 664504 186228 664556
rect 186280 664544 186286 664556
rect 197998 664544 198004 664556
rect 186280 664516 198004 664544
rect 186280 664504 186286 664516
rect 197998 664504 198004 664516
rect 198056 664504 198062 664556
rect 210234 664504 210240 664556
rect 210292 664544 210298 664556
rect 558914 664544 558920 664556
rect 210292 664516 558920 664544
rect 210292 664504 210298 664516
rect 558914 664504 558920 664516
rect 558972 664504 558978 664556
rect 9364 664448 175964 664476
rect 9364 664436 9370 664448
rect 180702 664436 180708 664488
rect 180760 664476 180766 664488
rect 534166 664476 534172 664488
rect 180760 664448 534172 664476
rect 180760 664436 180766 664448
rect 534166 664436 534172 664448
rect 534224 664436 534230 664488
rect 537386 664436 537392 664488
rect 537444 664476 537450 664488
rect 545114 664476 545120 664488
rect 537444 664448 545120 664476
rect 537444 664436 537450 664448
rect 545114 664436 545120 664448
rect 545172 664436 545178 664488
rect 6546 664368 6552 664420
rect 6604 664408 6610 664420
rect 195054 664408 195060 664420
rect 6604 664380 195060 664408
rect 6604 664368 6610 664380
rect 195054 664368 195060 664380
rect 195112 664368 195118 664420
rect 336734 664408 336740 664420
rect 316006 664380 336740 664408
rect 11698 664300 11704 664352
rect 11756 664340 11762 664352
rect 249518 664340 249524 664352
rect 11756 664312 249524 664340
rect 11756 664300 11762 664312
rect 249518 664300 249524 664312
rect 249576 664300 249582 664352
rect 264698 664300 264704 664352
rect 264756 664340 264762 664352
rect 316006 664340 316034 664380
rect 336734 664368 336740 664380
rect 336792 664368 336798 664420
rect 370682 664368 370688 664420
rect 370740 664408 370746 664420
rect 375374 664408 375380 664420
rect 370740 664380 375380 664408
rect 370740 664368 370746 664380
rect 375374 664368 375380 664380
rect 375432 664368 375438 664420
rect 376754 664368 376760 664420
rect 376812 664408 376818 664420
rect 391934 664408 391940 664420
rect 376812 664380 391940 664408
rect 376812 664368 376818 664380
rect 391934 664368 391940 664380
rect 391992 664368 391998 664420
rect 416130 664368 416136 664420
rect 416188 664408 416194 664420
rect 549990 664408 549996 664420
rect 416188 664380 549996 664408
rect 416188 664368 416194 664380
rect 549990 664368 549996 664380
rect 550048 664368 550054 664420
rect 264756 664312 316034 664340
rect 264756 664300 264762 664312
rect 349522 664300 349528 664352
rect 349580 664340 349586 664352
rect 548702 664340 548708 664352
rect 349580 664312 548708 664340
rect 349580 664300 349586 664312
rect 548702 664300 548708 664312
rect 548760 664300 548766 664352
rect 9398 664232 9404 664284
rect 9456 664272 9462 664284
rect 267734 664272 267740 664284
rect 9456 664244 267740 664272
rect 9456 664232 9462 664244
rect 267734 664232 267740 664244
rect 267792 664232 267798 664284
rect 322290 664232 322296 664284
rect 322348 664272 322354 664284
rect 551830 664272 551836 664284
rect 322348 664244 551836 664272
rect 322348 664232 322354 664244
rect 551830 664232 551836 664244
rect 551888 664232 551894 664284
rect 4982 664164 4988 664216
rect 5040 664204 5046 664216
rect 288894 664204 288900 664216
rect 5040 664176 288900 664204
rect 5040 664164 5046 664176
rect 288894 664164 288900 664176
rect 288952 664164 288958 664216
rect 291930 664164 291936 664216
rect 291988 664204 291994 664216
rect 551554 664204 551560 664216
rect 291988 664176 551560 664204
rect 291988 664164 291994 664176
rect 551554 664164 551560 664176
rect 551612 664164 551618 664216
rect 7650 664096 7656 664148
rect 7708 664136 7714 664148
rect 313274 664136 313280 664148
rect 7708 664108 313280 664136
rect 7708 664096 7714 664108
rect 313274 664096 313280 664108
rect 313332 664096 313338 664148
rect 319346 664096 319352 664148
rect 319404 664136 319410 664148
rect 549254 664136 549260 664148
rect 319404 664108 549260 664136
rect 319404 664096 319410 664108
rect 549254 664096 549260 664108
rect 549312 664096 549318 664148
rect 4798 664028 4804 664080
rect 4856 664068 4862 664080
rect 222289 664071 222347 664077
rect 222289 664068 222301 664071
rect 4856 664040 222301 664068
rect 4856 664028 4862 664040
rect 222289 664037 222301 664040
rect 222335 664037 222347 664071
rect 222289 664031 222347 664037
rect 222378 664028 222384 664080
rect 222436 664068 222442 664080
rect 552842 664068 552848 664080
rect 222436 664040 552848 664068
rect 222436 664028 222442 664040
rect 552842 664028 552848 664040
rect 552900 664028 552906 664080
rect 10410 663960 10416 664012
rect 10468 664000 10474 664012
rect 204070 664000 204076 664012
rect 10468 663972 204076 664000
rect 10468 663960 10474 663972
rect 204070 663960 204076 663972
rect 204128 663960 204134 664012
rect 213178 663960 213184 664012
rect 213236 664000 213242 664012
rect 548794 664000 548800 664012
rect 213236 663972 548800 664000
rect 213236 663960 213242 663972
rect 548794 663960 548800 663972
rect 548852 663960 548858 664012
rect 3418 663892 3424 663944
rect 3476 663932 3482 663944
rect 10502 663932 10508 663944
rect 3476 663904 10508 663932
rect 3476 663892 3482 663904
rect 10502 663892 10508 663904
rect 10560 663892 10566 663944
rect 10686 663892 10692 663944
rect 10744 663932 10750 663944
rect 382734 663932 382740 663944
rect 10744 663904 382740 663932
rect 10744 663892 10750 663904
rect 382734 663892 382740 663904
rect 382792 663892 382798 663944
rect 382829 663935 382887 663941
rect 382829 663901 382841 663935
rect 382875 663932 382887 663935
rect 548978 663932 548984 663944
rect 382875 663904 548984 663932
rect 382875 663901 382887 663904
rect 382829 663895 382887 663901
rect 548978 663892 548984 663904
rect 549036 663892 549042 663944
rect 4706 663824 4712 663876
rect 4764 663864 4770 663876
rect 131390 663864 131396 663876
rect 4764 663836 131396 663864
rect 4764 663824 4770 663836
rect 131390 663824 131396 663836
rect 131448 663824 131454 663876
rect 173802 663824 173808 663876
rect 173860 663864 173866 663876
rect 494790 663864 494796 663876
rect 173860 663836 382780 663864
rect 173860 663824 173866 663836
rect 38470 663756 38476 663808
rect 38528 663796 38534 663808
rect 43622 663796 43628 663808
rect 38528 663768 43628 663796
rect 38528 663756 38534 663768
rect 43622 663756 43628 663768
rect 43680 663756 43686 663808
rect 142154 663756 142160 663808
rect 142212 663796 142218 663808
rect 152550 663796 152556 663808
rect 142212 663768 152556 663796
rect 142212 663756 142218 663768
rect 152550 663756 152556 663768
rect 152608 663756 152614 663808
rect 222289 663799 222347 663805
rect 222289 663765 222301 663799
rect 222335 663796 222347 663799
rect 228358 663796 228364 663808
rect 222335 663768 228364 663796
rect 222335 663765 222347 663768
rect 222289 663759 222347 663765
rect 228358 663756 228364 663768
rect 228416 663756 228422 663808
rect 364794 663756 364800 663808
rect 364852 663796 364858 663808
rect 382645 663799 382703 663805
rect 382645 663796 382657 663799
rect 364852 663768 382657 663796
rect 364852 663756 364858 663768
rect 382645 663765 382657 663768
rect 382691 663765 382703 663799
rect 382752 663796 382780 663836
rect 383626 663836 494796 663864
rect 383626 663796 383654 663836
rect 494790 663824 494796 663836
rect 494848 663824 494854 663876
rect 507026 663824 507032 663876
rect 507084 663864 507090 663876
rect 550266 663864 550272 663876
rect 507084 663836 550272 663864
rect 507084 663824 507090 663836
rect 550266 663824 550272 663836
rect 550324 663824 550330 663876
rect 382752 663768 383654 663796
rect 382645 663759 382703 663765
rect 488810 663756 488816 663808
rect 488868 663796 488874 663808
rect 491294 663796 491300 663808
rect 488868 663768 491300 663796
rect 488868 663756 488874 663768
rect 491294 663756 491300 663768
rect 491352 663756 491358 663808
rect 540330 663756 540336 663808
rect 540388 663796 540394 663808
rect 542446 663796 542452 663808
rect 540388 663768 542452 663796
rect 540388 663756 540394 663768
rect 542446 663756 542452 663768
rect 542504 663756 542510 663808
rect 336734 663688 336740 663740
rect 336792 663728 336798 663740
rect 353294 663728 353300 663740
rect 336792 663700 353300 663728
rect 336792 663688 336798 663700
rect 353294 663688 353300 663700
rect 353352 663688 353358 663740
rect 355962 663688 355968 663740
rect 356020 663728 356026 663740
rect 546862 663728 546868 663740
rect 356020 663700 546868 663728
rect 356020 663688 356026 663700
rect 546862 663688 546868 663700
rect 546920 663688 546926 663740
rect 260742 663620 260748 663672
rect 260800 663660 260806 663672
rect 542722 663660 542728 663672
rect 260800 663632 542728 663660
rect 260800 663620 260806 663632
rect 542722 663620 542728 663632
rect 542780 663620 542786 663672
rect 261754 663552 261760 663604
rect 261812 663592 261818 663604
rect 580442 663592 580448 663604
rect 261812 663564 580448 663592
rect 261812 663552 261818 663564
rect 580442 663552 580448 663564
rect 580500 663552 580506 663604
rect 5258 663484 5264 663536
rect 5316 663524 5322 663536
rect 328270 663524 328276 663536
rect 5316 663496 328276 663524
rect 5316 663484 5322 663496
rect 328270 663484 328276 663496
rect 328328 663484 328334 663536
rect 339402 663484 339408 663536
rect 339460 663524 339466 663536
rect 543366 663524 543372 663536
rect 339460 663496 543372 663524
rect 339460 663484 339466 663496
rect 543366 663484 543372 663496
rect 543424 663484 543430 663536
rect 122466 663456 122472 663468
rect 122427 663428 122472 663456
rect 122466 663416 122472 663428
rect 122524 663416 122530 663468
rect 213822 663416 213828 663468
rect 213880 663456 213886 663468
rect 546678 663456 546684 663468
rect 213880 663428 546684 663456
rect 213880 663416 213886 663428
rect 546678 663416 546684 663428
rect 546736 663416 546742 663468
rect 39298 663348 39304 663400
rect 39356 663388 39362 663400
rect 372614 663388 372620 663400
rect 39356 663360 372620 663388
rect 39356 663348 39362 663360
rect 372614 663348 372620 663360
rect 372672 663348 372678 663400
rect 59262 663280 59268 663332
rect 59320 663320 59326 663332
rect 142154 663320 142160 663332
rect 59320 663292 142160 663320
rect 59320 663280 59326 663292
rect 142154 663280 142160 663292
rect 142212 663280 142218 663332
rect 209682 663280 209688 663332
rect 209740 663320 209746 663332
rect 545390 663320 545396 663332
rect 209740 663292 545396 663320
rect 209740 663280 209746 663292
rect 545390 663280 545396 663292
rect 545448 663280 545454 663332
rect 41138 663212 41144 663264
rect 41196 663252 41202 663264
rect 378134 663252 378140 663264
rect 41196 663224 378140 663252
rect 41196 663212 41202 663224
rect 378134 663212 378140 663224
rect 378192 663212 378198 663264
rect 40126 663144 40132 663196
rect 40184 663184 40190 663196
rect 434714 663184 434720 663196
rect 40184 663156 434720 663184
rect 40184 663144 40190 663156
rect 434714 663144 434720 663156
rect 434772 663144 434778 663196
rect 77202 663076 77208 663128
rect 77260 663116 77266 663128
rect 544010 663116 544016 663128
rect 77260 663088 544016 663116
rect 77260 663076 77266 663088
rect 544010 663076 544016 663088
rect 544068 663076 544074 663128
rect 53650 663008 53656 663060
rect 53708 663048 53714 663060
rect 546494 663048 546500 663060
rect 53708 663020 546500 663048
rect 53708 663008 53714 663020
rect 546494 663008 546500 663020
rect 546552 663008 546558 663060
rect 9490 662940 9496 662992
rect 9548 662980 9554 662992
rect 403710 662980 403716 662992
rect 9548 662952 403716 662980
rect 9548 662940 9554 662952
rect 403710 662940 403716 662952
rect 403768 662940 403774 662992
rect 5442 662872 5448 662924
rect 5500 662912 5506 662924
rect 409874 662912 409880 662924
rect 5500 662884 409880 662912
rect 5500 662872 5506 662884
rect 409874 662872 409880 662884
rect 409932 662872 409938 662924
rect 5350 662804 5356 662856
rect 5408 662844 5414 662856
rect 418798 662844 418804 662856
rect 5408 662816 418804 662844
rect 5408 662804 5414 662816
rect 418798 662804 418804 662816
rect 418856 662804 418862 662856
rect 433886 662844 433892 662856
rect 433847 662816 433892 662844
rect 433886 662804 433892 662816
rect 433944 662804 433950 662856
rect 479334 662844 479340 662856
rect 479295 662816 479340 662844
rect 479334 662804 479340 662816
rect 479392 662804 479398 662856
rect 95142 662736 95148 662788
rect 95200 662776 95206 662788
rect 547138 662776 547144 662788
rect 95200 662748 547144 662776
rect 95200 662736 95206 662748
rect 547138 662736 547144 662748
rect 547196 662736 547202 662788
rect 77202 662708 77208 662720
rect 77163 662680 77208 662708
rect 77202 662668 77208 662680
rect 77260 662668 77266 662720
rect 110414 662708 110420 662720
rect 110375 662680 110420 662708
rect 110414 662668 110420 662680
rect 110472 662668 110478 662720
rect 116762 662668 116768 662720
rect 116820 662708 116826 662720
rect 580350 662708 580356 662720
rect 116820 662680 580356 662708
rect 116820 662668 116826 662680
rect 580350 662668 580356 662680
rect 580408 662668 580414 662720
rect 49878 662640 49884 662652
rect 49839 662612 49884 662640
rect 49878 662600 49884 662612
rect 49936 662600 49942 662652
rect 59906 662640 59912 662652
rect 59867 662612 59912 662640
rect 59906 662600 59912 662612
rect 59964 662600 59970 662652
rect 68186 662600 68192 662652
rect 68244 662640 68250 662652
rect 548610 662640 548616 662652
rect 68244 662612 548616 662640
rect 68244 662600 68250 662612
rect 548610 662600 548616 662612
rect 548668 662600 548674 662652
rect 9122 662532 9128 662584
rect 9180 662572 9186 662584
rect 497550 662572 497556 662584
rect 9180 662544 497556 662572
rect 9180 662532 9186 662544
rect 497550 662532 497556 662544
rect 497608 662532 497614 662584
rect 506382 662572 506388 662584
rect 506343 662544 506388 662572
rect 506382 662532 506388 662544
rect 506440 662532 506446 662584
rect 543458 662504 543464 662516
rect 41386 662476 543464 662504
rect 40586 662328 40592 662380
rect 40644 662368 40650 662380
rect 41386 662368 41414 662476
rect 543458 662464 543464 662476
rect 543516 662464 543522 662516
rect 42705 662439 42763 662445
rect 42705 662405 42717 662439
rect 42751 662436 42763 662439
rect 544102 662436 544108 662448
rect 42751 662408 544108 662436
rect 42751 662405 42763 662408
rect 42705 662399 42763 662405
rect 544102 662396 544108 662408
rect 544160 662396 544166 662448
rect 40644 662340 41414 662368
rect 41601 662371 41659 662377
rect 40644 662328 40650 662340
rect 41601 662337 41613 662371
rect 41647 662368 41659 662371
rect 125594 662368 125600 662380
rect 41647 662340 125600 662368
rect 41647 662337 41659 662340
rect 41601 662331 41659 662337
rect 125594 662328 125600 662340
rect 125652 662328 125658 662380
rect 153841 662371 153899 662377
rect 153841 662337 153853 662371
rect 153887 662368 153899 662371
rect 155954 662368 155960 662380
rect 153887 662340 155960 662368
rect 153887 662337 153899 662340
rect 153841 662331 153899 662337
rect 155954 662328 155960 662340
rect 156012 662328 156018 662380
rect 354030 662368 354036 662380
rect 353991 662340 354036 662368
rect 354030 662328 354036 662340
rect 354088 662328 354094 662380
rect 358262 662368 358268 662380
rect 358223 662340 358268 662368
rect 358262 662328 358268 662340
rect 358320 662328 358326 662380
rect 425054 662368 425060 662380
rect 425015 662340 425060 662368
rect 425054 662328 425060 662340
rect 425112 662328 425118 662380
rect 426342 662328 426348 662380
rect 426400 662368 426406 662380
rect 546770 662368 546776 662380
rect 426400 662340 546776 662368
rect 426400 662328 426406 662340
rect 546770 662328 546776 662340
rect 546828 662328 546834 662380
rect 38930 662260 38936 662312
rect 38988 662300 38994 662312
rect 241514 662300 241520 662312
rect 38988 662272 241520 662300
rect 38988 662260 38994 662272
rect 241514 662260 241520 662272
rect 241572 662260 241578 662312
rect 310422 662260 310428 662312
rect 310480 662300 310486 662312
rect 545666 662300 545672 662312
rect 310480 662272 545672 662300
rect 310480 662260 310486 662272
rect 545666 662260 545672 662272
rect 545724 662260 545730 662312
rect 40678 662192 40684 662244
rect 40736 662232 40742 662244
rect 153841 662235 153899 662241
rect 153841 662232 153853 662235
rect 40736 662204 153853 662232
rect 40736 662192 40742 662204
rect 153841 662201 153853 662204
rect 153887 662201 153899 662235
rect 153841 662195 153899 662201
rect 155221 662235 155279 662241
rect 155221 662201 155233 662235
rect 155267 662232 155279 662235
rect 158530 662232 158536 662244
rect 155267 662204 158536 662232
rect 155267 662201 155279 662204
rect 155221 662195 155279 662201
rect 158530 662192 158536 662204
rect 158588 662192 158594 662244
rect 220722 662192 220728 662244
rect 220780 662232 220786 662244
rect 542630 662232 542636 662244
rect 220780 662204 542636 662232
rect 220780 662192 220786 662204
rect 542630 662192 542636 662204
rect 542688 662192 542694 662244
rect 40494 662124 40500 662176
rect 40552 662164 40558 662176
rect 245746 662164 245752 662176
rect 40552 662136 245752 662164
rect 40552 662124 40558 662136
rect 245746 662124 245752 662136
rect 245804 662124 245810 662176
rect 286410 662124 286416 662176
rect 286468 662164 286474 662176
rect 545758 662164 545764 662176
rect 286468 662136 545764 662164
rect 286468 662124 286474 662136
rect 545758 662124 545764 662136
rect 545816 662124 545822 662176
rect 8110 662056 8116 662108
rect 8168 662096 8174 662108
rect 128354 662096 128360 662108
rect 8168 662068 128360 662096
rect 8168 662056 8174 662068
rect 128354 662056 128360 662068
rect 128412 662056 128418 662108
rect 155862 662096 155868 662108
rect 155823 662068 155868 662096
rect 155862 662056 155868 662068
rect 155920 662056 155926 662108
rect 200022 662056 200028 662108
rect 200080 662096 200086 662108
rect 545482 662096 545488 662108
rect 200080 662068 545488 662096
rect 200080 662056 200086 662068
rect 545482 662056 545488 662068
rect 545540 662056 545546 662108
rect 7834 661988 7840 662040
rect 7892 662028 7898 662040
rect 309686 662028 309692 662040
rect 7892 662000 309692 662028
rect 7892 661988 7898 662000
rect 309686 661988 309692 662000
rect 309744 661988 309750 662040
rect 346946 661988 346952 662040
rect 347004 662028 347010 662040
rect 545206 662028 545212 662040
rect 347004 662000 545212 662028
rect 347004 661988 347010 662000
rect 545206 661988 545212 662000
rect 545264 661988 545270 662040
rect 6638 661920 6644 661972
rect 6696 661960 6702 661972
rect 200758 661960 200764 661972
rect 6696 661932 200764 661960
rect 6696 661920 6702 661932
rect 200758 661920 200764 661932
rect 200816 661920 200822 661972
rect 216582 661920 216588 661972
rect 216640 661960 216646 661972
rect 580258 661960 580264 661972
rect 216640 661932 580264 661960
rect 216640 661920 216646 661932
rect 580258 661920 580264 661932
rect 580316 661920 580322 661972
rect 37826 661852 37832 661904
rect 37884 661892 37890 661904
rect 471974 661892 471980 661904
rect 37884 661864 471980 661892
rect 37884 661852 37890 661864
rect 471974 661852 471980 661864
rect 472032 661852 472038 661904
rect 476022 661852 476028 661904
rect 476080 661892 476086 661904
rect 545942 661892 545948 661904
rect 476080 661864 545948 661892
rect 476080 661852 476086 661864
rect 545942 661852 545948 661864
rect 546000 661852 546006 661904
rect 4890 661784 4896 661836
rect 4948 661824 4954 661836
rect 379514 661824 379520 661836
rect 4948 661796 379520 661824
rect 4948 661784 4954 661796
rect 379514 661784 379520 661796
rect 379572 661784 379578 661836
rect 392394 661784 392400 661836
rect 392452 661824 392458 661836
rect 547322 661824 547328 661836
rect 392452 661796 547328 661824
rect 392452 661784 392458 661796
rect 547322 661784 547328 661796
rect 547380 661784 547386 661836
rect 4062 661716 4068 661768
rect 4120 661756 4126 661768
rect 400582 661756 400588 661768
rect 4120 661728 400588 661756
rect 4120 661716 4126 661728
rect 400582 661716 400588 661728
rect 400640 661716 400646 661768
rect 412542 661716 412548 661768
rect 412600 661756 412606 661768
rect 545574 661756 545580 661768
rect 412600 661728 545580 661756
rect 412600 661716 412606 661728
rect 545574 661716 545580 661728
rect 545632 661716 545638 661768
rect 37550 661648 37556 661700
rect 37608 661688 37614 661700
rect 511994 661688 512000 661700
rect 37608 661660 512000 661688
rect 37608 661648 37614 661660
rect 511994 661648 512000 661660
rect 512052 661648 512058 661700
rect 515214 661688 515220 661700
rect 515175 661660 515220 661688
rect 515214 661648 515220 661660
rect 515272 661648 515278 661700
rect 520182 661688 520188 661700
rect 520143 661660 520188 661688
rect 520182 661648 520188 661660
rect 520240 661648 520246 661700
rect 539594 661648 539600 661700
rect 539652 661688 539658 661700
rect 580718 661688 580724 661700
rect 539652 661660 580724 661688
rect 539652 661648 539658 661660
rect 580718 661648 580724 661660
rect 580776 661648 580782 661700
rect 3234 661580 3240 661632
rect 3292 661620 3298 661632
rect 425057 661623 425115 661629
rect 425057 661620 425069 661623
rect 3292 661592 425069 661620
rect 3292 661580 3298 661592
rect 425057 661589 425069 661592
rect 425103 661589 425115 661623
rect 425057 661583 425115 661589
rect 506385 661623 506443 661629
rect 506385 661589 506397 661623
rect 506431 661620 506443 661623
rect 543274 661620 543280 661632
rect 506431 661592 543280 661620
rect 506431 661589 506443 661592
rect 506385 661583 506443 661589
rect 543274 661580 543280 661592
rect 543332 661580 543338 661632
rect 6362 661512 6368 661564
rect 6420 661552 6426 661564
rect 155221 661555 155279 661561
rect 155221 661552 155233 661555
rect 6420 661524 155233 661552
rect 6420 661512 6426 661524
rect 155221 661521 155233 661524
rect 155267 661521 155279 661555
rect 155221 661515 155279 661521
rect 155865 661555 155923 661561
rect 155865 661521 155877 661555
rect 155911 661552 155923 661555
rect 427633 661555 427691 661561
rect 427633 661552 427645 661555
rect 155911 661524 427645 661552
rect 155911 661521 155923 661524
rect 155865 661515 155923 661521
rect 427633 661521 427645 661524
rect 427679 661521 427691 661555
rect 427633 661515 427691 661521
rect 427909 661555 427967 661561
rect 427909 661521 427921 661555
rect 427955 661552 427967 661555
rect 580534 661552 580540 661564
rect 427955 661524 580540 661552
rect 427955 661521 427967 661524
rect 427909 661515 427967 661521
rect 580534 661512 580540 661524
rect 580592 661512 580598 661564
rect 3970 661444 3976 661496
rect 4028 661484 4034 661496
rect 433889 661487 433947 661493
rect 433889 661484 433901 661487
rect 4028 661456 433901 661484
rect 4028 661444 4034 661456
rect 433889 661453 433901 661456
rect 433935 661453 433947 661487
rect 433889 661447 433947 661453
rect 520185 661487 520243 661493
rect 520185 661453 520197 661487
rect 520231 661484 520243 661487
rect 543090 661484 543096 661496
rect 520231 661456 543096 661484
rect 520231 661453 520243 661456
rect 520185 661447 520243 661453
rect 543090 661444 543096 661456
rect 543148 661444 543154 661496
rect 40218 661376 40224 661428
rect 40276 661416 40282 661428
rect 542998 661416 543004 661428
rect 40276 661388 543004 661416
rect 40276 661376 40282 661388
rect 542998 661376 543004 661388
rect 543056 661376 543062 661428
rect 41601 661351 41659 661357
rect 41601 661348 41613 661351
rect 41386 661320 41613 661348
rect 37366 661240 37372 661292
rect 37424 661280 37430 661292
rect 41386 661280 41414 661320
rect 41601 661317 41613 661320
rect 41647 661317 41659 661351
rect 41601 661311 41659 661317
rect 41690 661308 41696 661360
rect 41748 661348 41754 661360
rect 41748 661320 541296 661348
rect 41748 661308 41754 661320
rect 37424 661252 41414 661280
rect 42613 661283 42671 661289
rect 37424 661240 37430 661252
rect 42613 661249 42625 661283
rect 42659 661280 42671 661283
rect 541268 661280 541296 661320
rect 542262 661308 542268 661360
rect 542320 661348 542326 661360
rect 544378 661348 544384 661360
rect 542320 661320 544384 661348
rect 542320 661308 542326 661320
rect 544378 661308 544384 661320
rect 544436 661308 544442 661360
rect 544562 661280 544568 661292
rect 42659 661252 541204 661280
rect 541268 661252 544568 661280
rect 42659 661249 42671 661252
rect 42613 661243 42671 661249
rect 35894 661172 35900 661224
rect 35952 661212 35958 661224
rect 541069 661215 541127 661221
rect 541069 661212 541081 661215
rect 35952 661184 541081 661212
rect 35952 661172 35958 661184
rect 541069 661181 541081 661184
rect 541115 661181 541127 661215
rect 541069 661175 541127 661181
rect 3602 661104 3608 661156
rect 3660 661144 3666 661156
rect 479337 661147 479395 661153
rect 479337 661144 479349 661147
rect 3660 661116 479349 661144
rect 3660 661104 3666 661116
rect 479337 661113 479349 661116
rect 479383 661113 479395 661147
rect 541176 661144 541204 661252
rect 544562 661240 544568 661252
rect 544620 661240 544626 661292
rect 541253 661215 541311 661221
rect 541253 661181 541265 661215
rect 541299 661212 541311 661215
rect 542078 661212 542084 661224
rect 541299 661184 542084 661212
rect 541299 661181 541311 661184
rect 541253 661175 541311 661181
rect 542078 661172 542084 661184
rect 542136 661172 542142 661224
rect 544746 661144 544752 661156
rect 541176 661116 544752 661144
rect 479337 661107 479395 661113
rect 544746 661104 544752 661116
rect 544804 661104 544810 661156
rect 551462 661104 551468 661156
rect 551520 661144 551526 661156
rect 579614 661144 579620 661156
rect 551520 661116 579620 661144
rect 551520 661104 551526 661116
rect 579614 661104 579620 661116
rect 579672 661104 579678 661156
rect 39850 661036 39856 661088
rect 39908 661076 39914 661088
rect 41417 661079 41475 661085
rect 41417 661076 41429 661079
rect 39908 661048 41429 661076
rect 39908 661036 39914 661048
rect 41417 661045 41429 661048
rect 41463 661045 41475 661079
rect 41417 661039 41475 661045
rect 41877 661079 41935 661085
rect 41877 661045 41889 661079
rect 41923 661076 41935 661079
rect 49881 661079 49939 661085
rect 49881 661076 49893 661079
rect 41923 661048 49893 661076
rect 41923 661045 41935 661048
rect 41877 661039 41935 661045
rect 49881 661045 49893 661048
rect 49927 661045 49939 661079
rect 49881 661039 49939 661045
rect 77205 661079 77263 661085
rect 77205 661045 77217 661079
rect 77251 661076 77263 661079
rect 565814 661076 565820 661088
rect 77251 661048 565820 661076
rect 77251 661045 77263 661048
rect 77205 661039 77263 661045
rect 565814 661036 565820 661048
rect 565872 661036 565878 661088
rect 6822 660968 6828 661020
rect 6880 661008 6886 661020
rect 38746 661008 38752 661020
rect 6880 660980 38752 661008
rect 6880 660968 6886 660980
rect 38746 660968 38752 660980
rect 38804 660968 38810 661020
rect 41690 661008 41696 661020
rect 38856 660980 41696 661008
rect 37918 660900 37924 660952
rect 37976 660940 37982 660952
rect 38856 660940 38884 660980
rect 41690 660968 41696 660980
rect 41748 660968 41754 661020
rect 122469 661011 122527 661017
rect 122469 660977 122481 661011
rect 122515 661008 122527 661011
rect 515217 661011 515275 661017
rect 515217 661008 515229 661011
rect 122515 660980 515229 661008
rect 122515 660977 122527 660980
rect 122469 660971 122527 660977
rect 515217 660977 515229 660980
rect 515263 660977 515275 661011
rect 515217 660971 515275 660977
rect 37976 660912 38884 660940
rect 37976 660900 37982 660912
rect 40310 660900 40316 660952
rect 40368 660940 40374 660952
rect 53009 660943 53067 660949
rect 53009 660940 53021 660943
rect 40368 660912 53021 660940
rect 40368 660900 40374 660912
rect 53009 660909 53021 660912
rect 53055 660909 53067 660943
rect 53009 660903 53067 660909
rect 110417 660943 110475 660949
rect 110417 660909 110429 660943
rect 110463 660940 110475 660943
rect 354033 660943 354091 660949
rect 354033 660940 354045 660943
rect 110463 660912 354045 660940
rect 110463 660909 110475 660912
rect 110417 660903 110475 660909
rect 354033 660909 354045 660912
rect 354079 660909 354091 660943
rect 354033 660903 354091 660909
rect 37642 660832 37648 660884
rect 37700 660872 37706 660884
rect 46109 660875 46167 660881
rect 46109 660872 46121 660875
rect 37700 660844 46121 660872
rect 37700 660832 37706 660844
rect 46109 660841 46121 660844
rect 46155 660841 46167 660875
rect 46109 660835 46167 660841
rect 46201 660875 46259 660881
rect 46201 660841 46213 660875
rect 46247 660872 46259 660875
rect 59909 660875 59967 660881
rect 46247 660844 46704 660872
rect 46247 660841 46259 660844
rect 46201 660835 46259 660841
rect 39298 660804 39304 660816
rect 39259 660776 39304 660804
rect 39298 660764 39304 660776
rect 39356 660764 39362 660816
rect 41414 660764 41420 660816
rect 41472 660804 41478 660816
rect 46385 660807 46443 660813
rect 46385 660804 46397 660807
rect 41472 660776 46397 660804
rect 41472 660764 41478 660776
rect 46385 660773 46397 660776
rect 46431 660773 46443 660807
rect 46676 660804 46704 660844
rect 59909 660841 59921 660875
rect 59955 660872 59967 660875
rect 358265 660875 358323 660881
rect 358265 660872 358277 660875
rect 59955 660844 358277 660872
rect 59955 660841 59967 660844
rect 59909 660835 59967 660841
rect 358265 660841 358277 660844
rect 358311 660841 358323 660875
rect 541894 660872 541900 660884
rect 541855 660844 541900 660872
rect 358265 660835 358323 660841
rect 541894 660832 541900 660844
rect 541952 660832 541958 660884
rect 50893 660807 50951 660813
rect 50893 660804 50905 660807
rect 46676 660776 50905 660804
rect 46385 660767 46443 660773
rect 50893 660773 50905 660776
rect 50939 660773 50951 660807
rect 50893 660767 50951 660773
rect 51169 660807 51227 660813
rect 51169 660773 51181 660807
rect 51215 660804 51227 660807
rect 542262 660804 542268 660816
rect 51215 660776 542268 660804
rect 51215 660773 51227 660776
rect 51169 660767 51227 660773
rect 542262 660764 542268 660776
rect 542320 660764 542326 660816
rect 38194 660696 38200 660748
rect 38252 660736 38258 660748
rect 41509 660739 41567 660745
rect 38252 660708 41414 660736
rect 38252 660696 38258 660708
rect 41386 660668 41414 660708
rect 41509 660705 41521 660739
rect 41555 660736 41567 660739
rect 46201 660739 46259 660745
rect 46201 660736 46213 660739
rect 41555 660708 46213 660736
rect 41555 660705 41567 660708
rect 41509 660699 41567 660705
rect 46201 660705 46213 660708
rect 46247 660705 46259 660739
rect 46201 660699 46259 660705
rect 53009 660739 53067 660745
rect 53009 660705 53021 660739
rect 53055 660736 53067 660739
rect 541894 660736 541900 660748
rect 53055 660708 541900 660736
rect 53055 660705 53067 660708
rect 53009 660699 53067 660705
rect 541894 660696 541900 660708
rect 541952 660696 541958 660748
rect 46293 660671 46351 660677
rect 46293 660668 46305 660671
rect 41386 660640 46305 660668
rect 46293 660637 46305 660640
rect 46339 660637 46351 660671
rect 46293 660631 46351 660637
rect 46385 660671 46443 660677
rect 46385 660637 46397 660671
rect 46431 660668 46443 660671
rect 543550 660668 543556 660680
rect 46431 660640 543556 660668
rect 46431 660637 46443 660640
rect 46385 660631 46443 660637
rect 543550 660628 543556 660640
rect 543608 660628 543614 660680
rect 39298 660560 39304 660612
rect 39356 660600 39362 660612
rect 542538 660600 542544 660612
rect 39356 660572 542544 660600
rect 39356 660560 39362 660572
rect 542538 660560 542544 660572
rect 542596 660560 542602 660612
rect 40126 660492 40132 660544
rect 40184 660532 40190 660544
rect 40313 660535 40371 660541
rect 40313 660532 40325 660535
rect 40184 660504 40325 660532
rect 40184 660492 40190 660504
rect 40313 660501 40325 660504
rect 40359 660501 40371 660535
rect 40313 660495 40371 660501
rect 40770 660492 40776 660544
rect 40828 660532 40834 660544
rect 42705 660535 42763 660541
rect 42705 660532 42717 660535
rect 40828 660504 42717 660532
rect 40828 660492 40834 660504
rect 42705 660501 42717 660504
rect 42751 660501 42763 660535
rect 42705 660495 42763 660501
rect 46109 660535 46167 660541
rect 46109 660501 46121 660535
rect 46155 660532 46167 660535
rect 545298 660532 545304 660544
rect 46155 660504 545304 660532
rect 46155 660501 46167 660504
rect 46109 660495 46167 660501
rect 545298 660492 545304 660504
rect 545356 660492 545362 660544
rect 39022 660424 39028 660476
rect 39080 660464 39086 660476
rect 46201 660467 46259 660473
rect 46201 660464 46213 660467
rect 39080 660436 46213 660464
rect 39080 660424 39086 660436
rect 46201 660433 46213 660436
rect 46247 660433 46259 660467
rect 46201 660427 46259 660433
rect 46293 660467 46351 660473
rect 46293 660433 46305 660467
rect 46339 660464 46351 660467
rect 568574 660464 568580 660476
rect 46339 660436 568580 660464
rect 46339 660433 46351 660436
rect 46293 660427 46351 660433
rect 568574 660424 568580 660436
rect 568632 660424 568638 660476
rect 36998 660356 37004 660408
rect 37056 660396 37062 660408
rect 40586 660396 40592 660408
rect 37056 660368 40592 660396
rect 37056 660356 37062 660368
rect 40586 660356 40592 660368
rect 40644 660356 40650 660408
rect 40862 660356 40868 660408
rect 40920 660396 40926 660408
rect 580626 660396 580632 660408
rect 40920 660368 580632 660396
rect 40920 660356 40926 660368
rect 580626 660356 580632 660368
rect 580684 660356 580690 660408
rect 3878 660288 3884 660340
rect 3936 660328 3942 660340
rect 544930 660328 544936 660340
rect 3936 660300 544936 660328
rect 3936 660288 3942 660300
rect 544930 660288 544936 660300
rect 544988 660288 544994 660340
rect 37274 660220 37280 660272
rect 37332 660260 37338 660272
rect 42613 660263 42671 660269
rect 42613 660260 42625 660263
rect 37332 660232 42625 660260
rect 37332 660220 37338 660232
rect 42613 660229 42625 660232
rect 42659 660229 42671 660263
rect 42613 660223 42671 660229
rect 46201 660263 46259 660269
rect 46201 660229 46213 660263
rect 46247 660260 46259 660263
rect 542078 660260 542084 660272
rect 46247 660232 542084 660260
rect 46247 660229 46259 660232
rect 46201 660223 46259 660229
rect 542078 660220 542084 660232
rect 542136 660220 542142 660272
rect 542538 660220 542544 660272
rect 542596 660260 542602 660272
rect 542722 660260 542728 660272
rect 542596 660232 542728 660260
rect 542596 660220 542602 660232
rect 542722 660220 542728 660232
rect 542780 660220 542786 660272
rect 543369 660263 543427 660269
rect 543369 660229 543381 660263
rect 543415 660260 543427 660263
rect 543458 660260 543464 660272
rect 543415 660232 543464 660260
rect 543415 660229 543427 660232
rect 543369 660223 543427 660229
rect 543458 660220 543464 660232
rect 543516 660220 543522 660272
rect 39574 660152 39580 660204
rect 39632 660192 39638 660204
rect 543182 660192 543188 660204
rect 39632 660164 543188 660192
rect 39632 660152 39638 660164
rect 543182 660152 543188 660164
rect 543240 660152 543246 660204
rect 39114 660084 39120 660136
rect 39172 660124 39178 660136
rect 543458 660124 543464 660136
rect 39172 660096 543464 660124
rect 39172 660084 39178 660096
rect 543458 660084 543464 660096
rect 543516 660084 543522 660136
rect 544010 660084 544016 660136
rect 544068 660124 544074 660136
rect 544105 660127 544163 660133
rect 544105 660124 544117 660127
rect 544068 660096 544117 660124
rect 544068 660084 544074 660096
rect 544105 660093 544117 660096
rect 544151 660093 544163 660127
rect 544105 660087 544163 660093
rect 37734 660016 37740 660068
rect 37792 660056 37798 660068
rect 545022 660056 545028 660068
rect 37792 660028 545028 660056
rect 37792 660016 37798 660028
rect 545022 660016 545028 660028
rect 545080 660016 545086 660068
rect 39758 659948 39764 660000
rect 39816 659988 39822 660000
rect 549070 659988 549076 660000
rect 39816 659960 549076 659988
rect 39816 659948 39822 659960
rect 549070 659948 549076 659960
rect 549128 659948 549134 660000
rect 23474 659880 23480 659932
rect 23532 659920 23538 659932
rect 544470 659920 544476 659932
rect 23532 659892 544476 659920
rect 23532 659880 23538 659892
rect 544470 659880 544476 659892
rect 544528 659880 544534 659932
rect 6454 659812 6460 659864
rect 6512 659852 6518 659864
rect 544010 659852 544016 659864
rect 6512 659824 544016 659852
rect 6512 659812 6518 659824
rect 544010 659812 544016 659824
rect 544068 659812 544074 659864
rect 40126 659744 40132 659796
rect 40184 659784 40190 659796
rect 580166 659784 580172 659796
rect 40184 659756 580172 659784
rect 40184 659744 40190 659756
rect 580166 659744 580172 659756
rect 580224 659744 580230 659796
rect 3326 659676 3332 659728
rect 3384 659716 3390 659728
rect 546586 659716 546592 659728
rect 3384 659688 546592 659716
rect 3384 659676 3390 659688
rect 546586 659676 546592 659688
rect 546644 659676 546650 659728
rect 542722 659608 542728 659660
rect 542780 659648 542786 659660
rect 543366 659648 543372 659660
rect 542780 659620 543372 659648
rect 542780 659608 542786 659620
rect 543366 659608 543372 659620
rect 543424 659608 543430 659660
rect 544654 659608 544660 659660
rect 544712 659648 544718 659660
rect 580994 659648 581000 659660
rect 544712 659620 581000 659648
rect 544712 659608 544718 659620
rect 580994 659608 581000 659620
rect 581052 659608 581058 659660
rect 543366 659512 543372 659524
rect 543327 659484 543372 659512
rect 543366 659472 543372 659484
rect 543424 659472 543430 659524
rect 544102 659268 544108 659320
rect 544160 659308 544166 659320
rect 544746 659308 544752 659320
rect 544160 659280 544752 659308
rect 544160 659268 544166 659280
rect 544746 659268 544752 659280
rect 544804 659268 544810 659320
rect 544102 659172 544108 659184
rect 544063 659144 544108 659172
rect 544102 659132 544108 659144
rect 544160 659132 544166 659184
rect 40586 658656 40592 658708
rect 40644 658696 40650 658708
rect 41138 658696 41144 658708
rect 40644 658668 41144 658696
rect 40644 658656 40650 658668
rect 41138 658656 41144 658668
rect 41196 658656 41202 658708
rect 3418 658384 3424 658436
rect 3476 658424 3482 658436
rect 6730 658424 6736 658436
rect 3476 658396 6736 658424
rect 3476 658384 3482 658396
rect 6730 658384 6736 658396
rect 6788 658384 6794 658436
rect 38838 658384 38844 658436
rect 38896 658384 38902 658436
rect 36998 658288 37004 658300
rect 34440 658260 37004 658288
rect 32214 658180 32220 658232
rect 32272 658220 32278 658232
rect 34440 658220 34468 658260
rect 36998 658248 37004 658260
rect 37056 658248 37062 658300
rect 37734 658288 37740 658300
rect 37200 658260 37740 658288
rect 32272 658192 34468 658220
rect 32272 658180 32278 658192
rect 34514 658180 34520 658232
rect 34572 658220 34578 658232
rect 37200 658220 37228 658260
rect 37734 658248 37740 658260
rect 37792 658248 37798 658300
rect 34572 658192 37228 658220
rect 34572 658180 34578 658192
rect 37366 658112 37372 658164
rect 37424 658152 37430 658164
rect 37734 658152 37740 658164
rect 37424 658124 37740 658152
rect 37424 658112 37430 658124
rect 37734 658112 37740 658124
rect 37792 658112 37798 658164
rect 38856 658096 38884 658384
rect 38838 658044 38844 658096
rect 38896 658044 38902 658096
rect 41138 657364 41144 657416
rect 41196 657404 41202 657416
rect 41414 657404 41420 657416
rect 41196 657376 41420 657404
rect 41196 657364 41202 657376
rect 41414 657364 41420 657376
rect 41472 657364 41478 657416
rect 39298 657268 39304 657280
rect 39259 657240 39304 657268
rect 39298 657228 39304 657240
rect 39356 657228 39362 657280
rect 41414 657268 41420 657280
rect 41375 657240 41420 657268
rect 41414 657228 41420 657240
rect 41472 657228 41478 657280
rect 31018 657160 31024 657212
rect 31076 657200 31082 657212
rect 35802 657200 35808 657212
rect 31076 657172 35808 657200
rect 31076 657160 31082 657172
rect 35802 657160 35808 657172
rect 35860 657160 35866 657212
rect 38930 657160 38936 657212
rect 38988 657200 38994 657212
rect 40310 657200 40316 657212
rect 38988 657172 40316 657200
rect 38988 657160 38994 657172
rect 40310 657160 40316 657172
rect 40368 657160 40374 657212
rect 36906 657024 36912 657076
rect 36964 657064 36970 657076
rect 37274 657064 37280 657076
rect 36964 657036 37280 657064
rect 36964 657024 36970 657036
rect 37274 657024 37280 657036
rect 37332 657024 37338 657076
rect 40310 657064 40316 657076
rect 40271 657036 40316 657064
rect 40310 657024 40316 657036
rect 40368 657024 40374 657076
rect 19978 656888 19984 656940
rect 20036 656928 20042 656940
rect 23474 656928 23480 656940
rect 20036 656900 23480 656928
rect 20036 656888 20042 656900
rect 23474 656888 23480 656900
rect 23532 656888 23538 656940
rect 544102 655596 544108 655648
rect 544160 655636 544166 655648
rect 544565 655639 544623 655645
rect 544565 655636 544577 655639
rect 544160 655608 544577 655636
rect 544160 655596 544166 655608
rect 544565 655605 544577 655608
rect 544611 655605 544623 655639
rect 544565 655599 544623 655605
rect 32214 655568 32220 655580
rect 30392 655540 32220 655568
rect 29822 655460 29828 655512
rect 29880 655500 29886 655512
rect 30392 655500 30420 655540
rect 32214 655528 32220 655540
rect 32272 655528 32278 655580
rect 29880 655472 30420 655500
rect 29880 655460 29886 655472
rect 543642 655460 543648 655512
rect 543700 655500 543706 655512
rect 544102 655500 544108 655512
rect 543700 655472 544108 655500
rect 543700 655460 543706 655472
rect 544102 655460 544108 655472
rect 544160 655460 544166 655512
rect 38838 655324 38844 655376
rect 38896 655364 38902 655376
rect 40954 655364 40960 655376
rect 38896 655336 40960 655364
rect 38896 655324 38902 655336
rect 40954 655324 40960 655336
rect 41012 655324 41018 655376
rect 40770 655188 40776 655240
rect 40828 655228 40834 655240
rect 40954 655228 40960 655240
rect 40828 655200 40960 655228
rect 40828 655188 40834 655200
rect 40954 655188 40960 655200
rect 41012 655188 41018 655240
rect 544010 655052 544016 655104
rect 544068 655092 544074 655104
rect 544286 655092 544292 655104
rect 544068 655064 544292 655092
rect 544068 655052 544074 655064
rect 544286 655052 544292 655064
rect 544344 655052 544350 655104
rect 544286 654916 544292 654968
rect 544344 654956 544350 654968
rect 544562 654956 544568 654968
rect 544344 654928 544568 654956
rect 544344 654916 544350 654928
rect 544562 654916 544568 654928
rect 544620 654916 544626 654968
rect 544562 654820 544568 654832
rect 544523 654792 544568 654820
rect 544562 654780 544568 654792
rect 544620 654780 544626 654832
rect 33134 654576 33140 654628
rect 33192 654616 33198 654628
rect 34514 654616 34520 654628
rect 33192 654588 34520 654616
rect 33192 654576 33198 654588
rect 34514 654576 34520 654588
rect 34572 654576 34578 654628
rect 3418 654440 3424 654492
rect 3476 654480 3482 654492
rect 7558 654480 7564 654492
rect 3476 654452 7564 654480
rect 3476 654440 3482 654452
rect 7558 654440 7564 654452
rect 7616 654440 7622 654492
rect 3602 654412 3608 654424
rect 3436 654384 3608 654412
rect 3436 654356 3464 654384
rect 3602 654372 3608 654384
rect 3660 654372 3666 654424
rect 3418 654304 3424 654356
rect 3476 654304 3482 654356
rect 542170 654344 542176 654356
rect 542131 654316 542176 654344
rect 542170 654304 542176 654316
rect 542228 654304 542234 654356
rect 3234 654236 3240 654288
rect 3292 654276 3298 654288
rect 3602 654276 3608 654288
rect 3292 654248 3608 654276
rect 3292 654236 3298 654248
rect 3602 654236 3608 654248
rect 3660 654236 3666 654288
rect 541894 654236 541900 654288
rect 541952 654236 541958 654288
rect 32950 654168 32956 654220
rect 33008 654208 33014 654220
rect 36906 654208 36912 654220
rect 33008 654180 36912 654208
rect 33008 654168 33014 654180
rect 36906 654168 36912 654180
rect 36964 654168 36970 654220
rect 541912 654208 541940 654236
rect 541912 654180 542124 654208
rect 542096 654152 542124 654180
rect 41414 654140 41420 654152
rect 40788 654112 41420 654140
rect 40678 653964 40684 654016
rect 40736 654004 40742 654016
rect 40788 654004 40816 654112
rect 41414 654100 41420 654112
rect 41472 654100 41478 654152
rect 541897 654146 541955 654149
rect 541894 654094 541900 654146
rect 541952 654140 541958 654146
rect 541952 654106 541991 654140
rect 541952 654094 541958 654106
rect 542078 654100 542084 654152
rect 542136 654100 542142 654152
rect 40736 653976 40816 654004
rect 40736 653964 40742 653976
rect 37366 652740 37372 652792
rect 37424 652780 37430 652792
rect 38838 652780 38844 652792
rect 37424 652752 38844 652780
rect 37424 652740 37430 652752
rect 38838 652740 38844 652752
rect 38896 652740 38902 652792
rect 38933 652783 38991 652789
rect 38933 652749 38945 652783
rect 38979 652780 38991 652783
rect 40678 652780 40684 652792
rect 38979 652752 40684 652780
rect 38979 652749 38991 652752
rect 38933 652743 38991 652749
rect 40678 652740 40684 652752
rect 40736 652740 40742 652792
rect 17954 651380 17960 651432
rect 18012 651420 18018 651432
rect 19978 651420 19984 651432
rect 18012 651392 19984 651420
rect 18012 651380 18018 651392
rect 19978 651380 19984 651392
rect 20036 651380 20042 651432
rect 28994 651380 29000 651432
rect 29052 651420 29058 651432
rect 31018 651420 31024 651432
rect 29052 651392 31024 651420
rect 29052 651380 29058 651392
rect 31018 651380 31024 651392
rect 31076 651380 31082 651432
rect 562318 651380 562324 651432
rect 562376 651420 562382 651432
rect 562376 651392 564480 651420
rect 562376 651380 562382 651392
rect 3510 651312 3516 651364
rect 3568 651352 3574 651364
rect 38838 651352 38844 651364
rect 3568 651324 38844 651352
rect 3568 651312 3574 651324
rect 38838 651312 38844 651324
rect 38896 651312 38902 651364
rect 564452 651352 564480 651392
rect 567838 651352 567844 651364
rect 564452 651324 567844 651352
rect 567838 651312 567844 651324
rect 567896 651312 567902 651364
rect 542173 651287 542231 651293
rect 542173 651253 542185 651287
rect 542219 651284 542231 651287
rect 543642 651284 543648 651296
rect 542219 651256 543648 651284
rect 542219 651253 542231 651256
rect 542173 651247 542231 651253
rect 543642 651244 543648 651256
rect 543700 651244 543706 651296
rect 38838 650700 38844 650752
rect 38896 650740 38902 650752
rect 38933 650743 38991 650749
rect 38933 650740 38945 650743
rect 38896 650712 38945 650740
rect 38896 650700 38902 650712
rect 38933 650709 38945 650712
rect 38979 650709 38991 650743
rect 38933 650703 38991 650709
rect 26694 650020 26700 650072
rect 26752 650060 26758 650072
rect 29822 650060 29828 650072
rect 26752 650032 29828 650060
rect 26752 650020 26758 650032
rect 29822 650020 29828 650032
rect 29880 650020 29886 650072
rect 27062 648728 27068 648780
rect 27120 648768 27126 648780
rect 28994 648768 29000 648780
rect 27120 648740 29000 648768
rect 27120 648728 27126 648740
rect 28994 648728 29000 648740
rect 29052 648728 29058 648780
rect 567838 648592 567844 648644
rect 567896 648632 567902 648644
rect 567896 648604 568620 648632
rect 567896 648592 567902 648604
rect 36906 648524 36912 648576
rect 36964 648564 36970 648576
rect 37366 648564 37372 648576
rect 36964 648536 37372 648564
rect 36964 648524 36970 648536
rect 37366 648524 37372 648536
rect 37424 648524 37430 648576
rect 568592 648564 568620 648604
rect 571978 648564 571984 648576
rect 568592 648536 571984 648564
rect 571978 648524 571984 648536
rect 572036 648524 572042 648576
rect 37274 648456 37280 648508
rect 37332 648496 37338 648508
rect 38838 648496 38844 648508
rect 37332 648468 38844 648496
rect 37332 648456 37338 648468
rect 38838 648456 38844 648468
rect 38896 648456 38902 648508
rect 28258 647504 28264 647556
rect 28316 647544 28322 647556
rect 33134 647544 33140 647556
rect 28316 647516 33140 647544
rect 28316 647504 28322 647516
rect 33134 647504 33140 647516
rect 33192 647504 33198 647556
rect 31478 647232 31484 647284
rect 31536 647272 31542 647284
rect 32950 647272 32956 647284
rect 31536 647244 32956 647272
rect 31536 647232 31542 647244
rect 32950 647232 32956 647244
rect 33008 647232 33014 647284
rect 3694 647164 3700 647216
rect 3752 647204 3758 647216
rect 38838 647204 38844 647216
rect 3752 647176 38844 647204
rect 3752 647164 3758 647176
rect 38838 647164 38844 647176
rect 38896 647164 38902 647216
rect 24946 645940 24952 645992
rect 25004 645980 25010 645992
rect 27062 645980 27068 645992
rect 25004 645952 27068 645980
rect 25004 645940 25010 645952
rect 27062 645940 27068 645952
rect 27120 645940 27126 645992
rect 13814 645872 13820 645924
rect 13872 645912 13878 645924
rect 17862 645912 17868 645924
rect 13872 645884 17868 645912
rect 13872 645872 13878 645884
rect 17862 645872 17868 645884
rect 17920 645872 17926 645924
rect 26694 645912 26700 645924
rect 26206 645884 26700 645912
rect 22094 645804 22100 645856
rect 22152 645844 22158 645856
rect 26206 645844 26234 645884
rect 26694 645872 26700 645884
rect 26752 645872 26758 645924
rect 34514 645872 34520 645924
rect 34572 645912 34578 645924
rect 36906 645912 36912 645924
rect 34572 645884 36912 645912
rect 34572 645872 34578 645884
rect 36906 645872 36912 645884
rect 36964 645872 36970 645924
rect 22152 645816 26234 645844
rect 22152 645804 22158 645816
rect 29914 645192 29920 645244
rect 29972 645232 29978 645244
rect 31478 645232 31484 645244
rect 29972 645204 31484 645232
rect 29972 645192 29978 645204
rect 31478 645192 31484 645204
rect 31536 645192 31542 645244
rect 37366 643152 37372 643204
rect 37424 643192 37430 643204
rect 38838 643192 38844 643204
rect 37424 643164 38844 643192
rect 37424 643152 37430 643164
rect 38838 643152 38844 643164
rect 38896 643152 38902 643204
rect 30374 643084 30380 643136
rect 30432 643124 30438 643136
rect 34514 643124 34520 643136
rect 30432 643096 34520 643124
rect 30432 643084 30438 643096
rect 34514 643084 34520 643096
rect 34572 643084 34578 643136
rect 34606 643084 34612 643136
rect 34664 643124 34670 643136
rect 37274 643124 37280 643136
rect 34664 643096 37280 643124
rect 34664 643084 34670 643096
rect 37274 643084 37280 643096
rect 37332 643084 37338 643136
rect 3786 643016 3792 643068
rect 3844 643056 3850 643068
rect 38838 643056 38844 643068
rect 3844 643028 38844 643056
rect 3844 643016 3850 643028
rect 38838 643016 38844 643028
rect 38896 643016 38902 643068
rect 550082 641724 550088 641776
rect 550140 641764 550146 641776
rect 580074 641764 580080 641776
rect 550140 641736 580080 641764
rect 550140 641724 550146 641736
rect 580074 641724 580080 641736
rect 580132 641724 580138 641776
rect 27614 640364 27620 640416
rect 27672 640404 27678 640416
rect 30374 640404 30380 640416
rect 27672 640376 30380 640404
rect 27672 640364 27678 640376
rect 30374 640364 30380 640376
rect 30432 640364 30438 640416
rect 22738 640296 22744 640348
rect 22796 640336 22802 640348
rect 24946 640336 24952 640348
rect 22796 640308 24952 640336
rect 22796 640296 22802 640308
rect 24946 640296 24952 640308
rect 25004 640296 25010 640348
rect 28166 640296 28172 640348
rect 28224 640336 28230 640348
rect 29914 640336 29920 640348
rect 28224 640308 29920 640336
rect 28224 640296 28230 640308
rect 29914 640296 29920 640308
rect 29972 640296 29978 640348
rect 2774 640228 2780 640280
rect 2832 640268 2838 640280
rect 4890 640268 4896 640280
rect 2832 640240 4896 640268
rect 2832 640228 2838 640240
rect 4890 640228 4896 640240
rect 4948 640228 4954 640280
rect 11054 638936 11060 638988
rect 11112 638976 11118 638988
rect 13722 638976 13728 638988
rect 11112 638948 13728 638976
rect 11112 638936 11118 638948
rect 13722 638936 13728 638948
rect 13780 638936 13786 638988
rect 32950 638936 32956 638988
rect 33008 638976 33014 638988
rect 34606 638976 34612 638988
rect 33008 638948 34612 638976
rect 33008 638936 33014 638948
rect 34606 638936 34612 638948
rect 34664 638936 34670 638988
rect 11054 637616 11060 637628
rect 10336 637588 11060 637616
rect 8478 637508 8484 637560
rect 8536 637548 8542 637560
rect 10336 637548 10364 637588
rect 11054 637576 11060 637588
rect 11112 637576 11118 637628
rect 8536 637520 10364 637548
rect 8536 637508 8542 637520
rect 544838 637508 544844 637560
rect 544896 637548 544902 637560
rect 580902 637548 580908 637560
rect 544896 637520 580908 637548
rect 544896 637508 544902 637520
rect 580902 637508 580908 637520
rect 580960 637508 580966 637560
rect 20254 637304 20260 637356
rect 20312 637344 20318 637356
rect 22002 637344 22008 637356
rect 20312 637316 22008 637344
rect 20312 637304 20318 637316
rect 22002 637304 22008 637316
rect 22060 637304 22066 637356
rect 26234 637304 26240 637356
rect 26292 637344 26298 637356
rect 28166 637344 28172 637356
rect 26292 637316 28172 637344
rect 26292 637304 26298 637316
rect 28166 637304 28172 637316
rect 28224 637304 28230 637356
rect 37918 636256 37924 636268
rect 35866 636228 37924 636256
rect 35250 636148 35256 636200
rect 35308 636188 35314 636200
rect 35866 636188 35894 636228
rect 37918 636216 37924 636228
rect 37976 636216 37982 636268
rect 563698 636216 563704 636268
rect 563756 636256 563762 636268
rect 579982 636256 579988 636268
rect 563756 636228 579988 636256
rect 563756 636216 563762 636228
rect 579982 636216 579988 636228
rect 580040 636216 580046 636268
rect 35308 636160 35894 636188
rect 35308 636148 35314 636160
rect 30374 635128 30380 635180
rect 30432 635168 30438 635180
rect 32950 635168 32956 635180
rect 30432 635140 32956 635168
rect 30432 635128 30438 635140
rect 32950 635128 32956 635140
rect 33008 635128 33014 635180
rect 8478 634828 8484 634840
rect 7024 634800 8484 634828
rect 5534 634720 5540 634772
rect 5592 634760 5598 634772
rect 7024 634760 7052 634800
rect 8478 634788 8484 634800
rect 8536 634788 8542 634840
rect 27522 634828 27528 634840
rect 24872 634800 27528 634828
rect 5592 634732 7052 634760
rect 5592 634720 5598 634732
rect 23474 634720 23480 634772
rect 23532 634760 23538 634772
rect 24872 634760 24900 634800
rect 27522 634788 27528 634800
rect 27580 634788 27586 634840
rect 23532 634732 24900 634760
rect 23532 634720 23538 634732
rect 2774 633496 2780 633548
rect 2832 633536 2838 633548
rect 4890 633536 4896 633548
rect 2832 633508 4896 633536
rect 2832 633496 2838 633508
rect 4890 633496 4896 633508
rect 4948 633496 4954 633548
rect 35158 633468 35164 633480
rect 30392 633440 35164 633468
rect 30098 633360 30104 633412
rect 30156 633400 30162 633412
rect 30392 633400 30420 633440
rect 35158 633428 35164 633440
rect 35216 633428 35222 633480
rect 30156 633372 30420 633400
rect 30156 633360 30162 633372
rect 17218 632068 17224 632120
rect 17276 632108 17282 632120
rect 20254 632108 20260 632120
rect 17276 632080 20260 632108
rect 17276 632068 17282 632080
rect 20254 632068 20260 632080
rect 20312 632068 20318 632120
rect 23474 632108 23480 632120
rect 20732 632080 23480 632108
rect 19150 632000 19156 632052
rect 19208 632040 19214 632052
rect 20732 632040 20760 632080
rect 23474 632068 23480 632080
rect 23532 632068 23538 632120
rect 19208 632012 20760 632040
rect 19208 632000 19214 632012
rect 24854 631320 24860 631372
rect 24912 631360 24918 631372
rect 30282 631360 30288 631372
rect 24912 631332 30288 631360
rect 24912 631320 24918 631332
rect 30282 631320 30288 631332
rect 30340 631320 30346 631372
rect 26142 630680 26148 630692
rect 23860 630652 26148 630680
rect 3510 630572 3516 630624
rect 3568 630612 3574 630624
rect 7650 630612 7656 630624
rect 3568 630584 7656 630612
rect 3568 630572 3574 630584
rect 7650 630572 7656 630584
rect 7708 630572 7714 630624
rect 21358 630572 21364 630624
rect 21416 630612 21422 630624
rect 23860 630612 23888 630652
rect 26142 630640 26148 630652
rect 26200 630640 26206 630692
rect 26878 630640 26884 630692
rect 26936 630680 26942 630692
rect 30098 630680 30104 630692
rect 26936 630652 30104 630680
rect 26936 630640 26942 630652
rect 30098 630640 30104 630652
rect 30156 630640 30162 630692
rect 21416 630584 23888 630612
rect 21416 630572 21422 630584
rect 544102 629960 544108 630012
rect 544160 630000 544166 630012
rect 544838 630000 544844 630012
rect 544160 629972 544844 630000
rect 544160 629960 544166 629972
rect 544838 629960 544844 629972
rect 544896 629960 544902 630012
rect 4614 629892 4620 629944
rect 4672 629932 4678 629944
rect 5534 629932 5540 629944
rect 4672 629904 5540 629932
rect 4672 629892 4678 629904
rect 5534 629892 5540 629904
rect 5592 629892 5598 629944
rect 15838 629620 15844 629672
rect 15896 629660 15902 629672
rect 19150 629660 19156 629672
rect 15896 629632 19156 629660
rect 15896 629620 15902 629632
rect 19150 629620 19156 629632
rect 19208 629620 19214 629672
rect 571978 629212 571984 629264
rect 572036 629252 572042 629264
rect 575474 629252 575480 629264
rect 572036 629224 575480 629252
rect 572036 629212 572042 629224
rect 575474 629212 575480 629224
rect 575532 629212 575538 629264
rect 22094 627376 22100 627428
rect 22152 627416 22158 627428
rect 24762 627416 24768 627428
rect 22152 627388 24768 627416
rect 22152 627376 22158 627388
rect 24762 627376 24768 627388
rect 24820 627376 24826 627428
rect 575474 626560 575480 626612
rect 575532 626600 575538 626612
rect 576854 626600 576860 626612
rect 575532 626572 576860 626600
rect 575532 626560 575538 626572
rect 576854 626560 576860 626572
rect 576912 626560 576918 626612
rect 33778 626492 33784 626544
rect 33836 626532 33842 626544
rect 35250 626532 35256 626544
rect 33836 626504 35256 626532
rect 33836 626492 33842 626504
rect 35250 626492 35256 626504
rect 35308 626492 35314 626544
rect 32398 625200 32404 625252
rect 32456 625240 32462 625252
rect 37366 625240 37372 625252
rect 32456 625212 37372 625240
rect 32456 625200 32462 625212
rect 37366 625200 37372 625212
rect 37424 625200 37430 625252
rect 17954 623840 17960 623892
rect 18012 623880 18018 623892
rect 22738 623880 22744 623892
rect 18012 623852 22744 623880
rect 18012 623840 18018 623852
rect 22738 623840 22744 623852
rect 22796 623840 22802 623892
rect 19978 623772 19984 623824
rect 20036 623812 20042 623824
rect 22094 623812 22100 623824
rect 20036 623784 22100 623812
rect 20036 623772 20042 623784
rect 22094 623772 22100 623784
rect 22152 623772 22158 623824
rect 549070 623704 549076 623756
rect 549128 623744 549134 623756
rect 580166 623744 580172 623756
rect 549128 623716 580172 623744
rect 549128 623704 549134 623716
rect 580166 623704 580172 623716
rect 580224 623704 580230 623756
rect 15838 622452 15844 622464
rect 8312 622424 15844 622452
rect 8202 622344 8208 622396
rect 8260 622384 8266 622396
rect 8312 622384 8340 622424
rect 15838 622412 15844 622424
rect 15896 622412 15902 622464
rect 8260 622356 8340 622384
rect 8260 622344 8266 622356
rect 576854 621460 576860 621512
rect 576912 621500 576918 621512
rect 579522 621500 579528 621512
rect 576912 621472 579528 621500
rect 576912 621460 576918 621472
rect 579522 621460 579528 621472
rect 579580 621460 579586 621512
rect 20070 620984 20076 621036
rect 20128 621024 20134 621036
rect 21358 621024 21364 621036
rect 20128 620996 21364 621024
rect 20128 620984 20134 620996
rect 21358 620984 21364 620996
rect 21416 620984 21422 621036
rect 542262 620304 542268 620356
rect 542320 620344 542326 620356
rect 542630 620344 542636 620356
rect 542320 620316 542636 620344
rect 542320 620304 542326 620316
rect 542630 620304 542636 620316
rect 542688 620304 542694 620356
rect 15838 619556 15844 619608
rect 15896 619596 15902 619608
rect 17218 619596 17224 619608
rect 15896 619568 17224 619596
rect 15896 619556 15902 619568
rect 17218 619556 17224 619568
rect 17276 619556 17282 619608
rect 21358 619556 21364 619608
rect 21416 619596 21422 619608
rect 26878 619596 26884 619608
rect 21416 619568 26884 619596
rect 21416 619556 21422 619568
rect 26878 619556 26884 619568
rect 26936 619556 26942 619608
rect 3786 619488 3792 619540
rect 3844 619528 3850 619540
rect 8202 619528 8208 619540
rect 3844 619500 8208 619528
rect 3844 619488 3850 619500
rect 8202 619488 8208 619500
rect 8260 619488 8266 619540
rect 14458 619488 14464 619540
rect 14516 619528 14522 619540
rect 17862 619528 17868 619540
rect 14516 619500 17868 619528
rect 14516 619488 14522 619500
rect 17862 619488 17868 619500
rect 17920 619488 17926 619540
rect 25498 618264 25504 618316
rect 25556 618304 25562 618316
rect 38838 618304 38844 618316
rect 25556 618276 38844 618304
rect 25556 618264 25562 618276
rect 38838 618264 38844 618276
rect 38896 618264 38902 618316
rect 544838 618264 544844 618316
rect 544896 618304 544902 618316
rect 578878 618304 578884 618316
rect 544896 618276 578884 618304
rect 544896 618264 544902 618276
rect 578878 618264 578884 618276
rect 578936 618264 578942 618316
rect 3510 618196 3516 618248
rect 3568 618236 3574 618248
rect 4614 618236 4620 618248
rect 3568 618208 4620 618236
rect 3568 618196 3574 618208
rect 4614 618196 4620 618208
rect 4672 618196 4678 618248
rect 549898 616836 549904 616888
rect 549956 616876 549962 616888
rect 579982 616876 579988 616888
rect 549956 616848 579988 616876
rect 549956 616836 549962 616848
rect 579982 616836 579988 616848
rect 580040 616836 580046 616888
rect 3326 615408 3332 615460
rect 3384 615448 3390 615460
rect 32398 615448 32404 615460
rect 3384 615420 32404 615448
rect 3384 615408 3390 615420
rect 32398 615408 32404 615420
rect 32456 615408 32462 615460
rect 13814 614116 13820 614168
rect 13872 614156 13878 614168
rect 15838 614156 15844 614168
rect 13872 614128 15844 614156
rect 13872 614116 13878 614128
rect 15838 614116 15844 614128
rect 15896 614116 15902 614168
rect 18046 614116 18052 614168
rect 18104 614156 18110 614168
rect 20070 614156 20076 614168
rect 18104 614128 20076 614156
rect 18104 614116 18110 614128
rect 20070 614116 20076 614128
rect 20128 614116 20134 614168
rect 21358 614156 21364 614168
rect 20180 614128 21364 614156
rect 18782 614048 18788 614100
rect 18840 614088 18846 614100
rect 20180 614088 20208 614128
rect 21358 614116 21364 614128
rect 21416 614116 21422 614168
rect 22094 614116 22100 614168
rect 22152 614156 22158 614168
rect 28258 614156 28264 614168
rect 22152 614128 28264 614156
rect 22152 614116 22158 614128
rect 28258 614116 28264 614128
rect 28316 614116 28322 614168
rect 29638 614116 29644 614168
rect 29696 614156 29702 614168
rect 38838 614156 38844 614168
rect 29696 614128 38844 614156
rect 29696 614116 29702 614128
rect 38838 614116 38844 614128
rect 38896 614116 38902 614168
rect 18840 614060 20208 614088
rect 18840 614048 18846 614060
rect 546954 613368 546960 613420
rect 547012 613408 547018 613420
rect 580810 613408 580816 613420
rect 547012 613380 580816 613408
rect 547012 613368 547018 613380
rect 580810 613368 580816 613380
rect 580868 613368 580874 613420
rect 15838 611124 15844 611176
rect 15896 611164 15902 611176
rect 18046 611164 18052 611176
rect 15896 611136 18052 611164
rect 15896 611124 15902 611136
rect 18046 611124 18052 611136
rect 18104 611124 18110 611176
rect 3326 610104 3332 610156
rect 3384 610144 3390 610156
rect 8846 610144 8852 610156
rect 3384 610116 8852 610144
rect 3384 610104 3390 610116
rect 8846 610104 8852 610116
rect 8904 610104 8910 610156
rect 18782 610008 18788 610020
rect 16546 609980 18788 610008
rect 9030 609900 9036 609952
rect 9088 609940 9094 609952
rect 16546 609940 16574 609980
rect 18782 609968 18788 609980
rect 18840 609968 18846 610020
rect 9088 609912 16574 609940
rect 9088 609900 9094 609912
rect 11330 608200 11336 608252
rect 11388 608240 11394 608252
rect 13722 608240 13728 608252
rect 11388 608212 13728 608240
rect 11388 608200 11394 608212
rect 13722 608200 13728 608212
rect 13780 608200 13786 608252
rect 550358 607180 550364 607232
rect 550416 607220 550422 607232
rect 580166 607220 580172 607232
rect 550416 607192 580172 607220
rect 550416 607180 550422 607192
rect 580166 607180 580172 607192
rect 580224 607180 580230 607232
rect 17954 607112 17960 607164
rect 18012 607152 18018 607164
rect 19978 607152 19984 607164
rect 18012 607124 19984 607152
rect 18012 607112 18018 607124
rect 19978 607112 19984 607124
rect 20036 607112 20042 607164
rect 20162 606704 20168 606756
rect 20220 606744 20226 606756
rect 22002 606744 22008 606756
rect 20220 606716 22008 606744
rect 20220 606704 20226 606716
rect 22002 606704 22008 606716
rect 22060 606704 22066 606756
rect 544838 605956 544844 606008
rect 544896 605996 544902 606008
rect 546954 605996 546960 606008
rect 544896 605968 546960 605996
rect 544896 605956 544902 605968
rect 546954 605956 546960 605968
rect 547012 605956 547018 606008
rect 15194 605072 15200 605124
rect 15252 605112 15258 605124
rect 20162 605112 20168 605124
rect 15252 605084 20168 605112
rect 15252 605072 15258 605084
rect 20162 605072 20168 605084
rect 20220 605072 20226 605124
rect 13814 604596 13820 604648
rect 13872 604636 13878 604648
rect 17954 604636 17960 604648
rect 13872 604608 17960 604636
rect 13872 604596 13878 604608
rect 17954 604596 17960 604608
rect 18012 604596 18018 604648
rect 8202 604528 8208 604580
rect 8260 604568 8266 604580
rect 11330 604568 11336 604580
rect 8260 604540 11336 604568
rect 8260 604528 8266 604540
rect 11330 604528 11336 604540
rect 11388 604528 11394 604580
rect 13906 604528 13912 604580
rect 13964 604568 13970 604580
rect 15838 604568 15844 604580
rect 13964 604540 15844 604568
rect 13964 604528 13970 604540
rect 15838 604528 15844 604540
rect 15896 604528 15902 604580
rect 3326 604460 3332 604512
rect 3384 604500 3390 604512
rect 21358 604500 21364 604512
rect 3384 604472 21364 604500
rect 3384 604460 3390 604472
rect 21358 604460 21364 604472
rect 21416 604460 21422 604512
rect 548978 604392 548984 604444
rect 549036 604432 549042 604444
rect 579614 604432 579620 604444
rect 549036 604404 579620 604432
rect 549036 604392 549042 604404
rect 579614 604392 579620 604404
rect 579672 604392 579678 604444
rect 29730 603100 29736 603152
rect 29788 603140 29794 603152
rect 33778 603140 33784 603152
rect 29788 603112 33784 603140
rect 29788 603100 29794 603112
rect 33778 603100 33784 603112
rect 33836 603100 33842 603152
rect 11422 601740 11428 601792
rect 11480 601780 11486 601792
rect 13906 601780 13912 601792
rect 11480 601752 13912 601780
rect 11480 601740 11486 601752
rect 13906 601740 13912 601752
rect 13964 601740 13970 601792
rect 10962 601672 10968 601724
rect 11020 601712 11026 601724
rect 13814 601712 13820 601724
rect 11020 601684 13820 601712
rect 11020 601672 11026 601684
rect 13814 601672 13820 601684
rect 13872 601672 13878 601724
rect 3694 601604 3700 601656
rect 3752 601644 3758 601656
rect 38838 601644 38844 601656
rect 3752 601616 38844 601644
rect 3752 601604 3758 601616
rect 38838 601604 38844 601616
rect 38896 601604 38902 601656
rect 2774 601332 2780 601384
rect 2832 601372 2838 601384
rect 4706 601372 4712 601384
rect 2832 601344 4712 601372
rect 2832 601332 2838 601344
rect 4706 601332 4712 601344
rect 4764 601332 4770 601384
rect 543550 600924 543556 600976
rect 543608 600964 543614 600976
rect 558270 600964 558276 600976
rect 543608 600936 558276 600964
rect 543608 600924 543614 600936
rect 558270 600924 558276 600936
rect 558328 600924 558334 600976
rect 15194 600352 15200 600364
rect 13832 600324 15200 600352
rect 7650 600244 7656 600296
rect 7708 600284 7714 600296
rect 9030 600284 9036 600296
rect 7708 600256 9036 600284
rect 7708 600244 7714 600256
rect 9030 600244 9036 600256
rect 9088 600244 9094 600296
rect 13078 600244 13084 600296
rect 13136 600284 13142 600296
rect 13832 600284 13860 600324
rect 15194 600312 15200 600324
rect 15252 600312 15258 600364
rect 13136 600256 13860 600284
rect 13136 600244 13142 600256
rect 5534 597524 5540 597576
rect 5592 597564 5598 597576
rect 8202 597564 8208 597576
rect 5592 597536 8208 597564
rect 5592 597524 5598 597536
rect 8202 597524 8208 597536
rect 8260 597524 8266 597576
rect 558178 597524 558184 597576
rect 558236 597564 558242 597576
rect 580166 597564 580172 597576
rect 558236 597536 580172 597564
rect 558236 597524 558242 597536
rect 580166 597524 580172 597536
rect 580224 597524 580230 597576
rect 6730 597456 6736 597508
rect 6788 597496 6794 597508
rect 38838 597496 38844 597508
rect 6788 597468 38844 597496
rect 6788 597456 6794 597468
rect 38838 597456 38844 597468
rect 38896 597456 38902 597508
rect 558270 597456 558276 597508
rect 558328 597496 558334 597508
rect 562962 597496 562968 597508
rect 558328 597468 562968 597496
rect 558328 597456 558334 597468
rect 562962 597456 562968 597468
rect 563020 597456 563026 597508
rect 543642 596980 543648 597032
rect 543700 597020 543706 597032
rect 550082 597020 550088 597032
rect 543700 596992 550088 597020
rect 543700 596980 543706 596992
rect 550082 596980 550088 596992
rect 550140 596980 550146 597032
rect 10778 596776 10784 596828
rect 10836 596816 10842 596828
rect 11422 596816 11428 596828
rect 10836 596788 11428 596816
rect 10836 596776 10842 596788
rect 11422 596776 11428 596788
rect 11480 596776 11486 596828
rect 3326 595008 3332 595060
rect 3384 595048 3390 595060
rect 9214 595048 9220 595060
rect 3384 595020 9220 595048
rect 3384 595008 3390 595020
rect 9214 595008 9220 595020
rect 9272 595008 9278 595060
rect 10226 594804 10232 594856
rect 10284 594844 10290 594856
rect 13078 594844 13084 594856
rect 10284 594816 13084 594844
rect 10284 594804 10290 594816
rect 13078 594804 13084 594816
rect 13136 594804 13142 594856
rect 3326 593376 3332 593428
rect 3384 593416 3390 593428
rect 5534 593416 5540 593428
rect 3384 593388 5540 593416
rect 3384 593376 3390 593388
rect 5534 593376 5540 593388
rect 5592 593376 5598 593428
rect 562962 593308 562968 593360
rect 563020 593348 563026 593360
rect 579614 593348 579620 593360
rect 563020 593320 579620 593348
rect 563020 593308 563026 593320
rect 579614 593308 579620 593320
rect 579672 593308 579678 593360
rect 33778 592016 33784 592068
rect 33836 592056 33842 592068
rect 38838 592056 38844 592068
rect 33836 592028 38844 592056
rect 33836 592016 33842 592028
rect 38838 592016 38844 592028
rect 38896 592016 38902 592068
rect 8294 591064 8300 591116
rect 8352 591104 8358 591116
rect 10226 591104 10232 591116
rect 8352 591076 10232 591104
rect 8352 591064 8358 591076
rect 10226 591064 10232 591076
rect 10284 591064 10290 591116
rect 10962 590696 10968 590708
rect 8312 590668 10968 590696
rect 8018 590588 8024 590640
rect 8076 590628 8082 590640
rect 8312 590628 8340 590668
rect 10962 590656 10968 590668
rect 11020 590656 11026 590708
rect 8076 590600 8340 590628
rect 8076 590588 8082 590600
rect 3142 590316 3148 590368
rect 3200 590356 3206 590368
rect 6546 590356 6552 590368
rect 3200 590328 6552 590356
rect 3200 590316 3206 590328
rect 6546 590316 6552 590328
rect 6604 590316 6610 590368
rect 3878 589228 3884 589280
rect 3936 589268 3942 589280
rect 38838 589268 38844 589280
rect 3936 589240 38844 589268
rect 3936 589228 3942 589240
rect 38838 589228 38844 589240
rect 38896 589228 38902 589280
rect 28258 587936 28264 587988
rect 28316 587976 28322 587988
rect 29730 587976 29736 587988
rect 28316 587948 29736 587976
rect 28316 587936 28322 587948
rect 29730 587936 29736 587948
rect 29788 587936 29794 587988
rect 548978 587868 548984 587920
rect 549036 587908 549042 587920
rect 580166 587908 580172 587920
rect 549036 587880 580172 587908
rect 549036 587868 549042 587880
rect 580166 587868 580172 587880
rect 580224 587868 580230 587920
rect 14458 586548 14464 586560
rect 11072 586520 14464 586548
rect 9674 586440 9680 586492
rect 9732 586480 9738 586492
rect 11072 586480 11100 586520
rect 14458 586508 14464 586520
rect 14516 586508 14522 586560
rect 9732 586452 11100 586480
rect 9732 586440 9738 586452
rect 2774 585760 2780 585812
rect 2832 585800 2838 585812
rect 4982 585800 4988 585812
rect 2832 585772 4988 585800
rect 2832 585760 2838 585772
rect 4982 585760 4988 585772
rect 5040 585760 5046 585812
rect 3234 585148 3240 585200
rect 3292 585188 3298 585200
rect 8202 585188 8208 585200
rect 3292 585160 8208 585188
rect 3292 585148 3298 585160
rect 8202 585148 8208 585160
rect 8260 585148 8266 585200
rect 9030 583720 9036 583772
rect 9088 583760 9094 583772
rect 9674 583760 9680 583772
rect 9088 583732 9680 583760
rect 9088 583720 9094 583732
rect 9674 583720 9680 583732
rect 9732 583720 9738 583772
rect 38930 582836 38936 582888
rect 38988 582876 38994 582888
rect 40678 582876 40684 582888
rect 38988 582848 40684 582876
rect 38988 582836 38994 582848
rect 40678 582836 40684 582848
rect 40736 582836 40742 582888
rect 8018 582400 8024 582412
rect 6886 582372 8024 582400
rect 4154 582292 4160 582344
rect 4212 582332 4218 582344
rect 6886 582332 6914 582372
rect 8018 582360 8024 582372
rect 8076 582360 8082 582412
rect 545850 582360 545856 582412
rect 545908 582400 545914 582412
rect 579982 582400 579988 582412
rect 545908 582372 579988 582400
rect 545908 582360 545914 582372
rect 579982 582360 579988 582372
rect 580040 582360 580046 582412
rect 4212 582304 6914 582332
rect 4212 582292 4218 582304
rect 7650 581040 7656 581052
rect 6886 581012 7656 581040
rect 4246 580932 4252 580984
rect 4304 580972 4310 580984
rect 6886 580972 6914 581012
rect 7650 581000 7656 581012
rect 7708 581000 7714 581052
rect 4304 580944 6914 580972
rect 4304 580932 4310 580944
rect 3694 579640 3700 579692
rect 3752 579680 3758 579692
rect 4154 579680 4160 579692
rect 3752 579652 4160 579680
rect 3752 579640 3758 579652
rect 4154 579640 4160 579652
rect 4212 579640 4218 579692
rect 548886 579572 548892 579624
rect 548944 579612 548950 579624
rect 579614 579612 579620 579624
rect 548944 579584 579620 579612
rect 548944 579572 548950 579584
rect 579614 579572 579620 579584
rect 579672 579572 579678 579624
rect 3234 578688 3240 578740
rect 3292 578728 3298 578740
rect 4246 578728 4252 578740
rect 3292 578700 4252 578728
rect 3292 578688 3298 578700
rect 4246 578688 4252 578700
rect 4304 578688 4310 578740
rect 545298 578212 545304 578264
rect 545356 578252 545362 578264
rect 567838 578252 567844 578264
rect 545356 578224 567844 578252
rect 545356 578212 545362 578224
rect 567838 578212 567844 578224
rect 567896 578212 567902 578264
rect 8294 577124 8300 577176
rect 8352 577164 8358 577176
rect 10778 577164 10784 577176
rect 8352 577136 10784 577164
rect 8352 577124 8358 577136
rect 10778 577124 10784 577136
rect 10836 577124 10842 577176
rect 26878 575492 26884 575544
rect 26936 575532 26942 575544
rect 28258 575532 28264 575544
rect 26936 575504 28264 575532
rect 26936 575492 26942 575504
rect 28258 575492 28264 575504
rect 28316 575492 28322 575544
rect 545022 574880 545028 574932
rect 545080 574880 545086 574932
rect 545040 574784 545068 574880
rect 544856 574756 545068 574784
rect 544856 574580 544884 574756
rect 544930 574676 544936 574728
rect 544988 574716 544994 574728
rect 550358 574716 550364 574728
rect 544988 574688 550364 574716
rect 544988 574676 544994 574688
rect 550358 574676 550364 574688
rect 550416 574676 550422 574728
rect 544930 574580 544936 574592
rect 544856 574552 544936 574580
rect 544930 574540 544936 574552
rect 544988 574540 544994 574592
rect 8018 574132 8024 574184
rect 8076 574172 8082 574184
rect 9030 574172 9036 574184
rect 8076 574144 9036 574172
rect 8076 574132 8082 574144
rect 9030 574132 9036 574144
rect 9088 574132 9094 574184
rect 4982 574064 4988 574116
rect 5040 574104 5046 574116
rect 38838 574104 38844 574116
rect 5040 574076 38844 574104
rect 5040 574064 5046 574076
rect 38838 574064 38844 574076
rect 38896 574064 38902 574116
rect 4706 573724 4712 573776
rect 4764 573764 4770 573776
rect 8294 573764 8300 573776
rect 4764 573736 8300 573764
rect 4764 573724 4770 573736
rect 8294 573724 8300 573736
rect 8352 573724 8358 573776
rect 547230 572704 547236 572756
rect 547288 572744 547294 572756
rect 580166 572744 580172 572756
rect 547288 572716 580172 572744
rect 547288 572704 547294 572716
rect 580166 572704 580172 572716
rect 580224 572704 580230 572756
rect 3050 570256 3056 570308
rect 3108 570296 3114 570308
rect 7650 570296 7656 570308
rect 3108 570268 7656 570296
rect 3108 570256 3114 570268
rect 7650 570256 7656 570268
rect 7708 570256 7714 570308
rect 39114 568964 39120 569016
rect 39172 569004 39178 569016
rect 41506 569004 41512 569016
rect 39172 568976 41512 569004
rect 39172 568964 39178 568976
rect 41506 568964 41512 568976
rect 41564 568964 41570 569016
rect 8018 568596 8024 568608
rect 6886 568568 8024 568596
rect 4338 568488 4344 568540
rect 4396 568528 4402 568540
rect 6886 568528 6914 568568
rect 8018 568556 8024 568568
rect 8076 568556 8082 568608
rect 25590 568556 25596 568608
rect 25648 568596 25654 568608
rect 26878 568596 26884 568608
rect 25648 568568 26884 568596
rect 25648 568556 25654 568568
rect 26878 568556 26884 568568
rect 26936 568556 26942 568608
rect 4396 568500 6914 568528
rect 4396 568488 4402 568500
rect 2774 565972 2780 566024
rect 2832 566012 2838 566024
rect 5442 566012 5448 566024
rect 2832 565984 5448 566012
rect 2832 565972 2838 565984
rect 5442 565972 5448 565984
rect 5500 565972 5506 566024
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 4338 565876 4344 565888
rect 3108 565848 4344 565876
rect 3108 565836 3114 565848
rect 4338 565836 4344 565848
rect 4396 565836 4402 565888
rect 544930 565768 544936 565820
rect 544988 565808 544994 565820
rect 580626 565808 580632 565820
rect 544988 565780 580632 565808
rect 544988 565768 544994 565780
rect 580626 565768 580632 565780
rect 580684 565768 580690 565820
rect 3878 564408 3884 564460
rect 3936 564448 3942 564460
rect 4706 564448 4712 564460
rect 3936 564420 4712 564448
rect 3936 564408 3942 564420
rect 4706 564408 4712 564420
rect 4764 564408 4770 564460
rect 39942 562300 39948 562352
rect 40000 562340 40006 562352
rect 40218 562340 40224 562352
rect 40000 562312 40224 562340
rect 40000 562300 40006 562312
rect 40218 562300 40224 562312
rect 40276 562300 40282 562352
rect 3142 561620 3148 561672
rect 3200 561660 3206 561672
rect 38654 561660 38660 561672
rect 3200 561632 38660 561660
rect 3200 561620 3206 561632
rect 38654 561620 38660 561632
rect 38712 561620 38718 561672
rect 3142 560260 3148 560312
rect 3200 560300 3206 560312
rect 14458 560300 14464 560312
rect 3200 560272 14464 560300
rect 3200 560260 3206 560272
rect 14458 560260 14464 560272
rect 14516 560260 14522 560312
rect 21726 559784 21732 559836
rect 21784 559824 21790 559836
rect 25590 559824 25596 559836
rect 21784 559796 25596 559824
rect 21784 559784 21790 559796
rect 25590 559784 25596 559796
rect 25648 559784 25654 559836
rect 548702 558832 548708 558884
rect 548760 558872 548766 558884
rect 580166 558872 580172 558884
rect 548760 558844 580172 558872
rect 548760 558832 548766 558844
rect 580166 558832 580172 558844
rect 580224 558832 580230 558884
rect 24118 556180 24124 556232
rect 24176 556220 24182 556232
rect 38654 556220 38660 556232
rect 24176 556192 38660 556220
rect 24176 556180 24182 556192
rect 38654 556180 38660 556192
rect 38712 556180 38718 556232
rect 3142 556112 3148 556164
rect 3200 556152 3206 556164
rect 21726 556152 21732 556164
rect 3200 556124 21732 556152
rect 3200 556112 3206 556124
rect 21726 556112 21732 556124
rect 21784 556112 21790 556164
rect 556798 553392 556804 553444
rect 556856 553432 556862 553444
rect 580166 553432 580172 553444
rect 556856 553404 580172 553432
rect 556856 553392 556862 553404
rect 580166 553392 580172 553404
rect 580224 553392 580230 553444
rect 544930 552100 544936 552152
rect 544988 552140 544994 552152
rect 548978 552140 548984 552152
rect 544988 552112 548984 552140
rect 544988 552100 544994 552112
rect 548978 552100 548984 552112
rect 549036 552100 549042 552152
rect 3142 550740 3148 550792
rect 3200 550780 3206 550792
rect 6546 550780 6552 550792
rect 3200 550752 6552 550780
rect 3200 550740 3206 550752
rect 6546 550740 6552 550752
rect 6604 550740 6610 550792
rect 39942 548972 39948 549024
rect 40000 549012 40006 549024
rect 41322 549012 41328 549024
rect 40000 548984 41328 549012
rect 40000 548972 40006 548984
rect 41322 548972 41328 548984
rect 41380 548972 41386 549024
rect 544654 547680 544660 547732
rect 544712 547720 544718 547732
rect 544930 547720 544936 547732
rect 544712 547692 544936 547720
rect 544712 547680 544718 547692
rect 544930 547680 544936 547692
rect 544988 547680 544994 547732
rect 543458 547136 543464 547188
rect 543516 547176 543522 547188
rect 546034 547176 546040 547188
rect 543516 547148 546040 547176
rect 543516 547136 543522 547148
rect 546034 547136 546040 547148
rect 546092 547136 546098 547188
rect 544654 546456 544660 546508
rect 544712 546496 544718 546508
rect 562318 546496 562324 546508
rect 544712 546468 562324 546496
rect 544712 546456 544718 546468
rect 562318 546456 562324 546468
rect 562376 546456 562382 546508
rect 542170 543192 542176 543244
rect 542228 543232 542234 543244
rect 543458 543232 543464 543244
rect 542228 543204 543464 543232
rect 542228 543192 542234 543204
rect 543458 543192 543464 543204
rect 543516 543192 543522 543244
rect 3142 540948 3148 541000
rect 3200 540988 3206 541000
rect 35158 540988 35164 541000
rect 3200 540960 35164 540988
rect 3200 540948 3206 540960
rect 35158 540948 35164 540960
rect 35216 540948 35222 541000
rect 7742 539520 7748 539572
rect 7800 539560 7806 539572
rect 38654 539560 38660 539572
rect 7800 539532 38660 539560
rect 7800 539520 7806 539532
rect 38654 539520 38660 539532
rect 38712 539520 38718 539572
rect 548702 538840 548708 538892
rect 548760 538880 548766 538892
rect 580074 538880 580080 538892
rect 548760 538852 580080 538880
rect 548760 538840 548766 538852
rect 580074 538840 580080 538852
rect 580132 538840 580138 538892
rect 559558 538228 559564 538280
rect 559616 538268 559622 538280
rect 580166 538268 580172 538280
rect 559616 538240 580172 538268
rect 559616 538228 559622 538240
rect 580166 538228 580172 538240
rect 580224 538228 580230 538280
rect 546034 537480 546040 537532
rect 546092 537520 546098 537532
rect 553394 537520 553400 537532
rect 546092 537492 553400 537520
rect 546092 537480 546098 537492
rect 553394 537480 553400 537492
rect 553452 537480 553458 537532
rect 544654 535372 544660 535424
rect 544712 535412 544718 535424
rect 554038 535412 554044 535424
rect 544712 535384 554044 535412
rect 544712 535372 544718 535384
rect 554038 535372 554044 535384
rect 554096 535372 554102 535424
rect 553394 533332 553400 533384
rect 553452 533372 553458 533384
rect 565078 533372 565084 533384
rect 553452 533344 565084 533372
rect 553452 533332 553458 533344
rect 565078 533332 565084 533344
rect 565136 533332 565142 533384
rect 2774 531224 2780 531276
rect 2832 531264 2838 531276
rect 5350 531264 5356 531276
rect 2832 531236 5356 531264
rect 2832 531224 2838 531236
rect 5350 531224 5356 531236
rect 5408 531224 5414 531276
rect 6730 529932 6736 529984
rect 6788 529972 6794 529984
rect 38654 529972 38660 529984
rect 6788 529944 38660 529972
rect 6788 529932 6794 529944
rect 38654 529932 38660 529944
rect 38712 529932 38718 529984
rect 550450 528572 550456 528624
rect 550508 528612 550514 528624
rect 580166 528612 580172 528624
rect 550508 528584 580172 528612
rect 550508 528572 550514 528584
rect 580166 528572 580172 528584
rect 580224 528572 580230 528624
rect 565078 527076 565084 527128
rect 565136 527116 565142 527128
rect 569034 527116 569040 527128
rect 565136 527088 569040 527116
rect 565136 527076 565142 527088
rect 569034 527076 569040 527088
rect 569092 527076 569098 527128
rect 21358 525716 21364 525768
rect 21416 525756 21422 525768
rect 38654 525756 38660 525768
rect 21416 525728 38660 525756
rect 21416 525716 21422 525728
rect 38654 525716 38660 525728
rect 38712 525716 38718 525768
rect 569034 522928 569040 522980
rect 569092 522968 569098 522980
rect 571978 522968 571984 522980
rect 569092 522940 571984 522968
rect 569092 522928 569098 522940
rect 571978 522928 571984 522940
rect 572036 522928 572042 522980
rect 577498 521160 577504 521212
rect 577556 521200 577562 521212
rect 579614 521200 579620 521212
rect 577556 521172 579620 521200
rect 577556 521160 577562 521172
rect 579614 521160 579620 521172
rect 579672 521160 579678 521212
rect 544654 520820 544660 520872
rect 544712 520860 544718 520872
rect 548702 520860 548708 520872
rect 544712 520832 548708 520860
rect 544712 520820 544718 520832
rect 548702 520820 548708 520832
rect 548760 520820 548766 520872
rect 3142 520276 3148 520328
rect 3200 520316 3206 520328
rect 21358 520316 21364 520328
rect 3200 520288 21364 520316
rect 3200 520276 3206 520288
rect 21358 520276 21364 520288
rect 21416 520276 21422 520328
rect 571978 518168 571984 518220
rect 572036 518208 572042 518220
rect 580166 518208 580172 518220
rect 572036 518180 580172 518208
rect 572036 518168 572042 518180
rect 580166 518168 580172 518180
rect 580224 518168 580230 518220
rect 3142 516672 3148 516724
rect 3200 516712 3206 516724
rect 3694 516712 3700 516724
rect 3200 516684 3700 516712
rect 3200 516672 3206 516684
rect 3694 516672 3700 516684
rect 3752 516672 3758 516724
rect 3694 516400 3700 516452
rect 3752 516440 3758 516452
rect 9030 516440 9036 516452
rect 3752 516412 9036 516440
rect 3752 516400 3758 516412
rect 9030 516400 9036 516412
rect 9088 516400 9094 516452
rect 545022 516128 545028 516180
rect 545080 516168 545086 516180
rect 546126 516168 546132 516180
rect 545080 516140 546132 516168
rect 545080 516128 545086 516140
rect 546126 516128 546132 516140
rect 546184 516128 546190 516180
rect 544654 511844 544660 511896
rect 544712 511884 544718 511896
rect 545942 511884 545948 511896
rect 544712 511856 545948 511884
rect 544712 511844 544718 511856
rect 545942 511844 545948 511856
rect 546000 511844 546006 511896
rect 574094 509260 574100 509312
rect 574152 509300 574158 509312
rect 577498 509300 577504 509312
rect 574152 509272 577504 509300
rect 574152 509260 574158 509272
rect 577498 509260 577504 509272
rect 577556 509260 577562 509312
rect 3602 507424 3608 507476
rect 3660 507424 3666 507476
rect 3620 507272 3648 507424
rect 3602 507220 3608 507272
rect 3660 507220 3666 507272
rect 3510 507152 3516 507204
rect 3568 507192 3574 507204
rect 7926 507192 7932 507204
rect 3568 507164 7932 507192
rect 3568 507152 3574 507164
rect 7926 507152 7932 507164
rect 7984 507152 7990 507204
rect 563790 507084 563796 507136
rect 563848 507124 563854 507136
rect 574094 507124 574100 507136
rect 563848 507096 574100 507124
rect 563848 507084 563854 507096
rect 574094 507084 574100 507096
rect 574152 507084 574158 507136
rect 544654 506472 544660 506524
rect 544712 506512 544718 506524
rect 554130 506512 554136 506524
rect 544712 506484 554136 506512
rect 544712 506472 544718 506484
rect 554130 506472 554136 506484
rect 554188 506472 554194 506524
rect 542078 505928 542084 505980
rect 542136 505968 542142 505980
rect 542630 505968 542636 505980
rect 542136 505940 542636 505968
rect 542136 505928 542142 505940
rect 542630 505928 542636 505940
rect 542688 505928 542694 505980
rect 548702 503684 548708 503736
rect 548760 503724 548766 503736
rect 579982 503724 579988 503736
rect 548760 503696 579988 503724
rect 548760 503684 548766 503696
rect 579982 503684 579988 503696
rect 580040 503684 580046 503736
rect 549346 501576 549352 501628
rect 549404 501616 549410 501628
rect 580534 501616 580540 501628
rect 549404 501588 580540 501616
rect 549404 501576 549410 501588
rect 580534 501576 580540 501588
rect 580592 501576 580598 501628
rect 548794 500896 548800 500948
rect 548852 500936 548858 500948
rect 579706 500936 579712 500948
rect 548852 500908 579712 500936
rect 548852 500896 548858 500908
rect 579706 500896 579712 500908
rect 579764 500896 579770 500948
rect 8846 499468 8852 499520
rect 8904 499508 8910 499520
rect 38746 499508 38752 499520
rect 8904 499480 38752 499508
rect 8904 499468 8910 499480
rect 38746 499468 38752 499480
rect 38804 499468 38810 499520
rect 545022 498176 545028 498228
rect 545080 498216 545086 498228
rect 547782 498216 547788 498228
rect 545080 498188 547788 498216
rect 545080 498176 545086 498188
rect 547782 498176 547788 498188
rect 547840 498176 547846 498228
rect 26878 494028 26884 494080
rect 26936 494068 26942 494080
rect 38746 494068 38752 494080
rect 26936 494040 38752 494068
rect 26936 494028 26942 494040
rect 38746 494028 38752 494040
rect 38804 494028 38810 494080
rect 551646 494028 551652 494080
rect 551704 494068 551710 494080
rect 579982 494068 579988 494080
rect 551704 494040 579988 494068
rect 551704 494028 551710 494040
rect 579982 494028 579988 494040
rect 580040 494028 580046 494080
rect 544654 493892 544660 493944
rect 544712 493932 544718 493944
rect 549346 493932 549352 493944
rect 544712 493904 549352 493932
rect 544712 493892 544718 493904
rect 549346 493892 549352 493904
rect 549404 493892 549410 493944
rect 558914 492328 558920 492380
rect 558972 492368 558978 492380
rect 563790 492368 563796 492380
rect 558972 492340 563796 492368
rect 558972 492328 558978 492340
rect 563790 492328 563796 492340
rect 563848 492328 563854 492380
rect 554038 489880 554044 489932
rect 554096 489920 554102 489932
rect 580166 489920 580172 489932
rect 554096 489892 580172 489920
rect 554096 489880 554102 489892
rect 580166 489880 580172 489892
rect 580224 489880 580230 489932
rect 544654 489540 544660 489592
rect 544712 489580 544718 489592
rect 545666 489580 545672 489592
rect 544712 489552 545672 489580
rect 544712 489540 544718 489552
rect 545666 489540 545672 489552
rect 545724 489540 545730 489592
rect 8018 488520 8024 488572
rect 8076 488560 8082 488572
rect 38746 488560 38752 488572
rect 8076 488532 38752 488560
rect 8076 488520 8082 488532
rect 38746 488520 38752 488532
rect 38804 488520 38810 488572
rect 550818 488520 550824 488572
rect 550876 488560 550882 488572
rect 558914 488560 558920 488572
rect 550876 488532 558920 488560
rect 550876 488520 550882 488532
rect 558914 488520 558920 488532
rect 558972 488520 558978 488572
rect 543366 485800 543372 485852
rect 543424 485840 543430 485852
rect 545022 485840 545028 485852
rect 543424 485812 545028 485840
rect 543424 485800 543430 485812
rect 545022 485800 545028 485812
rect 545080 485800 545086 485852
rect 3510 485732 3516 485784
rect 3568 485772 3574 485784
rect 38746 485772 38752 485784
rect 3568 485744 38752 485772
rect 3568 485732 3574 485744
rect 38746 485732 38752 485744
rect 38804 485732 38810 485784
rect 548794 484372 548800 484424
rect 548852 484412 548858 484424
rect 580166 484412 580172 484424
rect 548852 484384 580172 484412
rect 548852 484372 548858 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 547506 478864 547512 478916
rect 547564 478904 547570 478916
rect 579614 478904 579620 478916
rect 547564 478876 579620 478904
rect 547564 478864 547570 478876
rect 579614 478864 579620 478876
rect 579672 478864 579678 478916
rect 545942 474716 545948 474768
rect 546000 474756 546006 474768
rect 580166 474756 580172 474768
rect 546000 474728 580172 474756
rect 546000 474716 546006 474728
rect 580166 474716 580172 474728
rect 580224 474716 580230 474768
rect 3510 471996 3516 472048
rect 3568 472036 3574 472048
rect 10778 472036 10784 472048
rect 3568 472008 10784 472036
rect 3568 471996 3574 472008
rect 10778 471996 10784 472008
rect 10836 471996 10842 472048
rect 2958 471860 2964 471912
rect 3016 471900 3022 471912
rect 3510 471900 3516 471912
rect 3016 471872 3516 471900
rect 3016 471860 3022 471872
rect 3510 471860 3516 471872
rect 3568 471860 3574 471912
rect 552934 469208 552940 469260
rect 552992 469248 552998 469260
rect 579982 469248 579988 469260
rect 552992 469220 579988 469248
rect 552992 469208 552998 469220
rect 579982 469208 579988 469220
rect 580040 469208 580046 469260
rect 3142 467304 3148 467356
rect 3200 467344 3206 467356
rect 7742 467344 7748 467356
rect 3200 467316 7748 467344
rect 3200 467304 3206 467316
rect 7742 467304 7748 467316
rect 7800 467304 7806 467356
rect 544654 466420 544660 466472
rect 544712 466460 544718 466472
rect 561030 466460 561036 466472
rect 544712 466432 561036 466460
rect 544712 466420 544718 466432
rect 561030 466420 561036 466432
rect 561088 466420 561094 466472
rect 2958 463632 2964 463684
rect 3016 463672 3022 463684
rect 38746 463672 38752 463684
rect 3016 463644 38752 463672
rect 3016 463632 3022 463644
rect 38746 463632 38752 463644
rect 38804 463632 38810 463684
rect 544654 462612 544660 462664
rect 544712 462652 544718 462664
rect 548794 462652 548800 462664
rect 544712 462624 548800 462652
rect 544712 462612 544718 462624
rect 548794 462612 548800 462624
rect 548852 462612 548858 462664
rect 3142 462408 3148 462460
rect 3200 462448 3206 462460
rect 7926 462448 7932 462460
rect 3200 462420 7932 462448
rect 3200 462408 3206 462420
rect 7926 462408 7932 462420
rect 7984 462408 7990 462460
rect 547598 460844 547604 460896
rect 547656 460884 547662 460896
rect 580166 460884 580172 460896
rect 547656 460856 580172 460884
rect 547656 460844 547662 460856
rect 580166 460844 580172 460856
rect 580224 460844 580230 460896
rect 3050 459484 3056 459536
rect 3108 459524 3114 459536
rect 38746 459524 38752 459536
rect 3108 459496 38752 459524
rect 3108 459484 3114 459496
rect 38746 459484 38752 459496
rect 38804 459484 38810 459536
rect 543458 458804 543464 458856
rect 543516 458844 543522 458856
rect 562042 458844 562048 458856
rect 543516 458816 562048 458844
rect 543516 458804 543522 458816
rect 562042 458804 562048 458816
rect 562100 458804 562106 458856
rect 562042 455404 562048 455456
rect 562100 455444 562106 455456
rect 566458 455444 566464 455456
rect 562100 455416 566464 455444
rect 562100 455404 562106 455416
rect 566458 455404 566464 455416
rect 566516 455404 566522 455456
rect 39942 455336 39948 455388
rect 40000 455376 40006 455388
rect 41230 455376 41236 455388
rect 40000 455348 41236 455376
rect 40000 455336 40006 455348
rect 41230 455336 41236 455348
rect 41288 455336 41294 455388
rect 550082 454044 550088 454096
rect 550140 454084 550146 454096
rect 580166 454084 580172 454096
rect 550140 454056 580172 454084
rect 550140 454044 550146 454056
rect 580166 454044 580172 454056
rect 580224 454044 580230 454096
rect 3234 452888 3240 452940
rect 3292 452928 3298 452940
rect 9582 452928 9588 452940
rect 3292 452900 9588 452928
rect 3292 452888 3298 452900
rect 9582 452888 9588 452900
rect 9640 452888 9646 452940
rect 544654 452616 544660 452668
rect 544712 452656 544718 452668
rect 574738 452656 574744 452668
rect 544712 452628 574744 452656
rect 544712 452616 544718 452628
rect 574738 452616 574744 452628
rect 574796 452616 574802 452668
rect 548794 449896 548800 449948
rect 548852 449936 548858 449948
rect 580166 449936 580172 449948
rect 548852 449908 580172 449936
rect 548852 449896 548858 449908
rect 580166 449896 580172 449908
rect 580224 449896 580230 449948
rect 544654 449828 544660 449880
rect 544712 449868 544718 449880
rect 580534 449868 580540 449880
rect 544712 449840 580540 449868
rect 544712 449828 544718 449840
rect 580534 449828 580540 449840
rect 580592 449828 580598 449880
rect 37458 449216 37464 449268
rect 37516 449256 37522 449268
rect 39298 449256 39304 449268
rect 37516 449228 39304 449256
rect 37516 449216 37522 449228
rect 39298 449216 39304 449228
rect 39356 449216 39362 449268
rect 3142 447108 3148 447160
rect 3200 447148 3206 447160
rect 13078 447148 13084 447160
rect 3200 447120 13084 447148
rect 3200 447108 3206 447120
rect 13078 447108 13084 447120
rect 13136 447108 13142 447160
rect 3234 444388 3240 444440
rect 3292 444428 3298 444440
rect 38746 444428 38752 444440
rect 3292 444400 38752 444428
rect 3292 444388 3298 444400
rect 38746 444388 38752 444400
rect 38804 444388 38810 444440
rect 547598 444388 547604 444440
rect 547656 444428 547662 444440
rect 580166 444428 580172 444440
rect 547656 444400 580172 444428
rect 547656 444388 547662 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 566458 442212 566464 442264
rect 566516 442252 566522 442264
rect 574094 442252 574100 442264
rect 566516 442224 574100 442252
rect 566516 442212 566522 442224
rect 574094 442212 574100 442224
rect 574152 442212 574158 442264
rect 544930 440308 544936 440360
rect 544988 440348 544994 440360
rect 550082 440348 550088 440360
rect 544988 440320 550088 440348
rect 544988 440308 544994 440320
rect 550082 440308 550088 440320
rect 550140 440308 550146 440360
rect 39482 440240 39488 440292
rect 39540 440280 39546 440292
rect 41046 440280 41052 440292
rect 39540 440252 41052 440280
rect 39540 440240 39546 440252
rect 41046 440240 41052 440252
rect 41104 440240 41110 440292
rect 551738 440240 551744 440292
rect 551796 440280 551802 440292
rect 580166 440280 580172 440292
rect 551796 440252 580172 440280
rect 551796 440240 551802 440252
rect 580166 440240 580172 440252
rect 580224 440240 580230 440292
rect 3234 438812 3240 438864
rect 3292 438852 3298 438864
rect 11698 438852 11704 438864
rect 3292 438824 11704 438852
rect 3292 438812 3298 438824
rect 11698 438812 11704 438824
rect 11756 438812 11762 438864
rect 574094 437384 574100 437436
rect 574152 437424 574158 437436
rect 577498 437424 577504 437436
rect 574152 437396 577504 437424
rect 574152 437384 574158 437396
rect 577498 437384 577504 437396
rect 577556 437384 577562 437436
rect 543918 435684 543924 435736
rect 543976 435724 543982 435736
rect 545574 435724 545580 435736
rect 543976 435696 545580 435724
rect 543976 435684 543982 435696
rect 545574 435684 545580 435696
rect 545632 435684 545638 435736
rect 550082 434732 550088 434784
rect 550140 434772 550146 434784
rect 580166 434772 580172 434784
rect 550140 434744 580172 434772
rect 550140 434732 550146 434744
rect 580166 434732 580172 434744
rect 580224 434732 580230 434784
rect 2958 431876 2964 431928
rect 3016 431916 3022 431928
rect 38746 431916 38752 431928
rect 3016 431888 38752 431916
rect 3016 431876 3022 431888
rect 38746 431876 38752 431888
rect 38804 431876 38810 431928
rect 577498 431400 577504 431452
rect 577556 431440 577562 431452
rect 579614 431440 579620 431452
rect 577556 431412 579620 431440
rect 577556 431400 577562 431412
rect 579614 431400 579620 431412
rect 579672 431400 579678 431452
rect 543918 431332 543924 431384
rect 543976 431372 543982 431384
rect 545482 431372 545488 431384
rect 543976 431344 545488 431372
rect 543976 431332 543982 431344
rect 545482 431332 545488 431344
rect 545540 431332 545546 431384
rect 3234 429020 3240 429072
rect 3292 429060 3298 429072
rect 6730 429060 6736 429072
rect 3292 429032 6736 429060
rect 3292 429020 3298 429032
rect 6730 429020 6736 429032
rect 6788 429020 6794 429072
rect 21450 426436 21456 426488
rect 21508 426476 21514 426488
rect 38746 426476 38752 426488
rect 21508 426448 38752 426476
rect 21508 426436 21514 426448
rect 38746 426436 38752 426448
rect 38804 426436 38810 426488
rect 548886 425076 548892 425128
rect 548944 425116 548950 425128
rect 580166 425116 580172 425128
rect 548944 425088 580172 425116
rect 548944 425076 548950 425088
rect 580166 425076 580172 425088
rect 580224 425076 580230 425128
rect 3234 423308 3240 423360
rect 3292 423348 3298 423360
rect 9490 423348 9496 423360
rect 3292 423320 9496 423348
rect 3292 423308 3298 423320
rect 9490 423308 9496 423320
rect 9548 423308 9554 423360
rect 41046 418140 41052 418192
rect 41104 418180 41110 418192
rect 41690 418180 41696 418192
rect 41104 418152 41696 418180
rect 41104 418140 41110 418152
rect 41690 418140 41696 418152
rect 41748 418140 41754 418192
rect 3234 418072 3240 418124
rect 3292 418112 3298 418124
rect 9398 418112 9404 418124
rect 3292 418084 9404 418112
rect 3292 418072 3298 418084
rect 9398 418072 9404 418084
rect 9456 418072 9462 418124
rect 544194 417732 544200 417784
rect 544252 417772 544258 417784
rect 546862 417772 546868 417784
rect 544252 417744 546868 417772
rect 544252 417732 544258 417744
rect 546862 417732 546868 417744
rect 546920 417732 546926 417784
rect 3142 413652 3148 413704
rect 3200 413692 3206 413704
rect 6638 413692 6644 413704
rect 3200 413664 6644 413692
rect 3200 413652 3206 413664
rect 6638 413652 6644 413664
rect 6696 413652 6702 413704
rect 9582 412632 9588 412684
rect 9640 412672 9646 412684
rect 38746 412672 38752 412684
rect 9640 412644 38752 412672
rect 9640 412632 9646 412644
rect 38746 412632 38752 412644
rect 38804 412632 38810 412684
rect 552566 409844 552572 409896
rect 552624 409884 552630 409896
rect 580166 409884 580172 409896
rect 552624 409856 580172 409884
rect 552624 409844 552630 409856
rect 580166 409844 580172 409856
rect 580224 409844 580230 409896
rect 544194 409028 544200 409080
rect 544252 409068 544258 409080
rect 546770 409068 546776 409080
rect 544252 409040 546776 409068
rect 544252 409028 544258 409040
rect 546770 409028 546776 409040
rect 546828 409028 546834 409080
rect 2774 408348 2780 408400
rect 2832 408388 2838 408400
rect 5166 408388 5172 408400
rect 2832 408360 5172 408388
rect 2832 408348 2838 408360
rect 5166 408348 5172 408360
rect 5224 408348 5230 408400
rect 39390 405900 39396 405952
rect 39448 405940 39454 405952
rect 41138 405940 41144 405952
rect 39448 405912 41144 405940
rect 39448 405900 39454 405912
rect 41138 405900 41144 405912
rect 41196 405900 41202 405952
rect 553118 405696 553124 405748
rect 553176 405736 553182 405748
rect 580166 405736 580172 405748
rect 553176 405708 580172 405736
rect 553176 405696 553182 405708
rect 580166 405696 580172 405708
rect 580224 405696 580230 405748
rect 544930 405628 544936 405680
rect 544988 405668 544994 405680
rect 552566 405668 552572 405680
rect 544988 405640 552572 405668
rect 544988 405628 544994 405640
rect 552566 405628 552572 405640
rect 552624 405628 552630 405680
rect 3234 404268 3240 404320
rect 3292 404308 3298 404320
rect 29638 404308 29644 404320
rect 3292 404280 29644 404308
rect 3292 404268 3298 404280
rect 29638 404268 29644 404280
rect 29696 404268 29702 404320
rect 562318 401548 562324 401600
rect 562376 401588 562382 401600
rect 579706 401588 579712 401600
rect 562376 401560 579712 401588
rect 562376 401548 562382 401560
rect 579706 401548 579712 401560
rect 579764 401548 579770 401600
rect 544838 400392 544844 400444
rect 544896 400392 544902 400444
rect 544856 400240 544884 400392
rect 544838 400188 544844 400240
rect 544896 400188 544902 400240
rect 544746 400120 544752 400172
rect 544804 400160 544810 400172
rect 553118 400160 553124 400172
rect 544804 400132 553124 400160
rect 544804 400120 544810 400132
rect 553118 400120 553124 400132
rect 553176 400120 553182 400172
rect 6822 398828 6828 398880
rect 6880 398868 6886 398880
rect 38746 398868 38752 398880
rect 6880 398840 38752 398868
rect 6880 398828 6886 398840
rect 38746 398828 38752 398840
rect 38804 398828 38810 398880
rect 3234 398556 3240 398608
rect 3292 398596 3298 398608
rect 9306 398596 9312 398608
rect 3292 398568 9312 398596
rect 3292 398556 3298 398568
rect 9306 398556 9312 398568
rect 9364 398556 9370 398608
rect 569862 398080 569868 398132
rect 569920 398120 569926 398132
rect 580626 398120 580632 398132
rect 569920 398092 580632 398120
rect 569920 398080 569926 398092
rect 580626 398080 580632 398092
rect 580684 398080 580690 398132
rect 544930 397400 544936 397452
rect 544988 397440 544994 397452
rect 550358 397440 550364 397452
rect 544988 397412 550364 397440
rect 544988 397400 544994 397412
rect 550358 397400 550364 397412
rect 550416 397400 550422 397452
rect 544746 395972 544752 396024
rect 544804 396012 544810 396024
rect 551738 396012 551744 396024
rect 544804 395984 551744 396012
rect 544804 395972 544810 395984
rect 551738 395972 551744 395984
rect 551796 395972 551802 396024
rect 557534 395292 557540 395344
rect 557592 395332 557598 395344
rect 569862 395332 569868 395344
rect 557592 395304 569868 395332
rect 557592 395292 557598 395304
rect 569862 395292 569868 395304
rect 569920 395292 569926 395344
rect 2774 393592 2780 393644
rect 2832 393632 2838 393644
rect 5166 393632 5172 393644
rect 2832 393604 5172 393632
rect 2832 393592 2838 393604
rect 5166 393592 5172 393604
rect 5224 393592 5230 393644
rect 550358 391212 550364 391264
rect 550416 391252 550422 391264
rect 563054 391252 563060 391264
rect 550416 391224 563060 391252
rect 550416 391212 550422 391224
rect 563054 391212 563060 391224
rect 563112 391212 563118 391264
rect 551186 390804 551192 390856
rect 551244 390844 551250 390856
rect 557534 390844 557540 390856
rect 551244 390816 557540 390844
rect 551244 390804 551250 390816
rect 557534 390804 557540 390816
rect 557592 390804 557598 390856
rect 544746 390600 544752 390652
rect 544804 390640 544810 390652
rect 551922 390640 551928 390652
rect 544804 390612 551928 390640
rect 544804 390600 544810 390612
rect 551922 390600 551928 390612
rect 551980 390600 551986 390652
rect 551738 390532 551744 390584
rect 551796 390572 551802 390584
rect 579614 390572 579620 390584
rect 551796 390544 579620 390572
rect 551796 390532 551802 390544
rect 579614 390532 579620 390544
rect 579672 390532 579678 390584
rect 563054 388424 563060 388476
rect 563112 388464 563118 388476
rect 570598 388464 570604 388476
rect 563112 388436 570604 388464
rect 563112 388424 563118 388436
rect 570598 388424 570604 388436
rect 570656 388424 570662 388476
rect 548978 386384 548984 386436
rect 549036 386424 549042 386436
rect 580166 386424 580172 386436
rect 549036 386396 580172 386424
rect 549036 386384 549042 386396
rect 580166 386384 580172 386396
rect 580224 386384 580230 386436
rect 548334 386112 548340 386164
rect 548392 386152 548398 386164
rect 551186 386152 551192 386164
rect 548392 386124 551192 386152
rect 548392 386112 548398 386124
rect 551186 386112 551192 386124
rect 551244 386112 551250 386164
rect 2774 384752 2780 384804
rect 2832 384792 2838 384804
rect 5258 384792 5264 384804
rect 2832 384764 5264 384792
rect 2832 384752 2838 384764
rect 5258 384752 5264 384764
rect 5316 384752 5322 384804
rect 543182 382576 543188 382628
rect 543240 382616 543246 382628
rect 550542 382616 550548 382628
rect 543240 382588 550548 382616
rect 543240 382576 543246 382588
rect 550542 382576 550548 382588
rect 550600 382576 550606 382628
rect 570598 382168 570604 382220
rect 570656 382208 570662 382220
rect 579798 382208 579804 382220
rect 570656 382180 579804 382208
rect 570656 382168 570662 382180
rect 579798 382168 579804 382180
rect 579856 382168 579862 382220
rect 546034 380944 546040 380996
rect 546092 380984 546098 380996
rect 548334 380984 548340 380996
rect 546092 380956 548340 380984
rect 546092 380944 546098 380956
rect 548334 380944 548340 380956
rect 548392 380944 548398 380996
rect 550542 378088 550548 378140
rect 550600 378128 550606 378140
rect 552566 378128 552572 378140
rect 550600 378100 552572 378128
rect 550600 378088 550606 378100
rect 552566 378088 552572 378100
rect 552624 378088 552630 378140
rect 544746 377476 544752 377528
rect 544804 377516 544810 377528
rect 550174 377516 550180 377528
rect 544804 377488 550180 377516
rect 544804 377476 544810 377488
rect 550174 377476 550180 377488
rect 550232 377476 550238 377528
rect 550266 376660 550272 376712
rect 550324 376700 550330 376712
rect 580166 376700 580172 376712
rect 550324 376672 580172 376700
rect 550324 376660 550330 376672
rect 580166 376660 580172 376672
rect 580224 376660 580230 376712
rect 552566 374892 552572 374944
rect 552624 374932 552630 374944
rect 558362 374932 558368 374944
rect 552624 374904 558368 374932
rect 552624 374892 552630 374904
rect 558362 374892 558368 374904
rect 558420 374892 558426 374944
rect 551830 372512 551836 372564
rect 551888 372552 551894 372564
rect 579614 372552 579620 372564
rect 551888 372524 579620 372552
rect 551888 372512 551894 372524
rect 579614 372512 579620 372524
rect 579672 372512 579678 372564
rect 3234 368500 3240 368552
rect 3292 368540 3298 368552
rect 33870 368540 33876 368552
rect 3292 368512 33876 368540
rect 3292 368500 3298 368512
rect 33870 368500 33876 368512
rect 33928 368500 33934 368552
rect 551830 365712 551836 365764
rect 551888 365752 551894 365764
rect 580166 365752 580172 365764
rect 551888 365724 580172 365752
rect 551888 365712 551894 365724
rect 580166 365712 580172 365724
rect 580224 365712 580230 365764
rect 544746 364148 544752 364200
rect 544804 364188 544810 364200
rect 545390 364188 545396 364200
rect 544804 364160 545396 364188
rect 544804 364148 544810 364160
rect 545390 364148 545396 364160
rect 545448 364148 545454 364200
rect 544838 362924 544844 362976
rect 544896 362964 544902 362976
rect 545390 362964 545396 362976
rect 544896 362936 545396 362964
rect 544896 362924 544902 362936
rect 545390 362924 545396 362936
rect 545448 362924 545454 362976
rect 574830 361564 574836 361616
rect 574888 361604 574894 361616
rect 580166 361604 580172 361616
rect 574888 361576 580172 361604
rect 574888 361564 574894 361576
rect 580166 361564 580172 361576
rect 580224 361564 580230 361616
rect 544930 358776 544936 358828
rect 544988 358816 544994 358828
rect 560938 358816 560944 358828
rect 544988 358788 560944 358816
rect 544988 358776 544994 358788
rect 560938 358776 560944 358788
rect 560996 358776 561002 358828
rect 550174 356056 550180 356108
rect 550232 356096 550238 356108
rect 579982 356096 579988 356108
rect 550232 356068 579988 356096
rect 550232 356056 550238 356068
rect 579982 356056 579988 356068
rect 580040 356056 580046 356108
rect 3142 354628 3148 354680
rect 3200 354668 3206 354680
rect 10870 354668 10876 354680
rect 3200 354640 10876 354668
rect 3200 354628 3206 354640
rect 10870 354628 10876 354640
rect 10928 354628 10934 354680
rect 561030 353200 561036 353252
rect 561088 353240 561094 353252
rect 580166 353240 580172 353252
rect 561088 353212 580172 353240
rect 561088 353200 561094 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 558270 352520 558276 352572
rect 558328 352560 558334 352572
rect 574830 352560 574836 352572
rect 558328 352532 574836 352560
rect 558328 352520 558334 352532
rect 574830 352520 574836 352532
rect 574888 352520 574894 352572
rect 6638 350548 6644 350600
rect 6696 350588 6702 350600
rect 38746 350588 38752 350600
rect 6696 350560 38752 350588
rect 6696 350548 6702 350560
rect 38746 350548 38752 350560
rect 38804 350548 38810 350600
rect 558362 350140 558368 350192
rect 558420 350180 558426 350192
rect 561030 350180 561036 350192
rect 558420 350152 561036 350180
rect 558420 350140 558426 350152
rect 561030 350140 561036 350152
rect 561088 350140 561094 350192
rect 2774 349188 2780 349240
rect 2832 349228 2838 349240
rect 5258 349228 5264 349240
rect 2832 349200 5264 349228
rect 2832 349188 2838 349200
rect 5258 349188 5264 349200
rect 5316 349188 5322 349240
rect 5350 346400 5356 346452
rect 5408 346440 5414 346452
rect 38746 346440 38752 346452
rect 5408 346412 38752 346440
rect 5408 346400 5414 346412
rect 38746 346400 38752 346412
rect 38804 346400 38810 346452
rect 553302 346400 553308 346452
rect 553360 346440 553366 346452
rect 580166 346440 580172 346452
rect 553360 346412 580172 346440
rect 553360 346400 553366 346412
rect 580166 346400 580172 346412
rect 580224 346400 580230 346452
rect 3326 344360 3332 344412
rect 3384 344400 3390 344412
rect 9306 344400 9312 344412
rect 3384 344372 9312 344400
rect 3384 344360 3390 344372
rect 9306 344360 9312 344372
rect 9364 344360 9370 344412
rect 544746 342184 544752 342236
rect 544804 342224 544810 342236
rect 553302 342224 553308 342236
rect 544804 342196 553308 342224
rect 544804 342184 544810 342196
rect 553302 342184 553308 342196
rect 553360 342184 553366 342236
rect 561030 340824 561036 340876
rect 561088 340864 561094 340876
rect 569218 340864 569224 340876
rect 561088 340836 569224 340864
rect 561088 340824 561094 340836
rect 569218 340824 569224 340836
rect 569276 340824 569282 340876
rect 3326 339464 3332 339516
rect 3384 339504 3390 339516
rect 9398 339504 9404 339516
rect 3384 339476 9404 339504
rect 3384 339464 3390 339476
rect 9398 339464 9404 339476
rect 9456 339464 9462 339516
rect 546126 338036 546132 338088
rect 546184 338076 546190 338088
rect 580166 338076 580172 338088
rect 546184 338048 580172 338076
rect 546184 338036 546190 338048
rect 580166 338036 580172 338048
rect 580224 338036 580230 338088
rect 542998 336676 543004 336728
rect 543056 336716 543062 336728
rect 546402 336716 546408 336728
rect 543056 336688 546408 336716
rect 543056 336676 543062 336688
rect 546402 336676 546408 336688
rect 546460 336676 546466 336728
rect 2958 334840 2964 334892
rect 3016 334880 3022 334892
rect 6454 334880 6460 334892
rect 3016 334852 6460 334880
rect 3016 334840 3022 334852
rect 6454 334840 6460 334852
rect 6512 334840 6518 334892
rect 569218 334364 569224 334416
rect 569276 334404 569282 334416
rect 574094 334404 574100 334416
rect 569276 334376 574100 334404
rect 569276 334364 569282 334376
rect 574094 334364 574100 334376
rect 574152 334364 574158 334416
rect 3326 332596 3332 332648
rect 3384 332636 3390 332648
rect 38746 332636 38752 332648
rect 3384 332608 38752 332636
rect 3384 332596 3390 332608
rect 38746 332596 38752 332608
rect 38804 332596 38810 332648
rect 541894 330964 541900 331016
rect 541952 331004 541958 331016
rect 547690 331004 547696 331016
rect 541952 330976 547696 331004
rect 541952 330964 541958 330976
rect 547690 330964 547696 330976
rect 547748 330964 547754 331016
rect 39574 329740 39580 329792
rect 39632 329780 39638 329792
rect 40770 329780 40776 329792
rect 39632 329752 40776 329780
rect 39632 329740 39638 329752
rect 40770 329740 40776 329752
rect 40828 329740 40834 329792
rect 3234 328720 3240 328772
rect 3292 328760 3298 328772
rect 6454 328760 6460 328772
rect 3292 328732 6460 328760
rect 3292 328720 3298 328732
rect 6454 328720 6460 328732
rect 6512 328720 6518 328772
rect 574094 328380 574100 328432
rect 574152 328420 574158 328432
rect 579982 328420 579988 328432
rect 574152 328392 579988 328420
rect 574152 328380 574158 328392
rect 579982 328380 579988 328392
rect 580040 328380 580046 328432
rect 37090 324232 37096 324284
rect 37148 324272 37154 324284
rect 38746 324272 38752 324284
rect 37148 324244 38752 324272
rect 37148 324232 37154 324244
rect 38746 324232 38752 324244
rect 38804 324232 38810 324284
rect 547690 322872 547696 322924
rect 547748 322912 547754 322924
rect 579798 322912 579804 322924
rect 547748 322884 579804 322912
rect 547748 322872 547754 322884
rect 579798 322872 579804 322884
rect 579856 322872 579862 322924
rect 544930 318928 544936 318980
rect 544988 318968 544994 318980
rect 550266 318968 550272 318980
rect 544988 318940 550272 318968
rect 544988 318928 544994 318940
rect 550266 318928 550272 318940
rect 550324 318928 550330 318980
rect 37458 318792 37464 318844
rect 37516 318832 37522 318844
rect 39298 318832 39304 318844
rect 37516 318804 39304 318832
rect 37516 318792 37522 318804
rect 39298 318792 39304 318804
rect 39356 318792 39362 318844
rect 546126 316684 546132 316736
rect 546184 316724 546190 316736
rect 558270 316724 558276 316736
rect 546184 316696 558276 316724
rect 546184 316684 546190 316696
rect 558270 316684 558276 316696
rect 558328 316684 558334 316736
rect 3326 315936 3332 315988
rect 3384 315976 3390 315988
rect 26878 315976 26884 315988
rect 3384 315948 26884 315976
rect 3384 315936 3390 315948
rect 26878 315936 26884 315948
rect 26936 315936 26942 315988
rect 2958 314644 2964 314696
rect 3016 314684 3022 314696
rect 38746 314684 38752 314696
rect 3016 314656 38752 314684
rect 3016 314644 3022 314656
rect 38746 314644 38752 314656
rect 38804 314644 38810 314696
rect 575474 313896 575480 313948
rect 575532 313936 575538 313948
rect 580718 313936 580724 313948
rect 575532 313908 580724 313936
rect 575532 313896 575538 313908
rect 580718 313896 580724 313908
rect 580776 313896 580782 313948
rect 551922 313216 551928 313268
rect 551980 313256 551986 313268
rect 580166 313256 580172 313268
rect 551980 313228 580172 313256
rect 551980 313216 551986 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 559650 311108 559656 311160
rect 559708 311148 559714 311160
rect 575474 311148 575480 311160
rect 559708 311120 575480 311148
rect 559708 311108 559714 311120
rect 575474 311108 575480 311120
rect 575532 311108 575538 311160
rect 3326 310496 3332 310548
rect 3384 310536 3390 310548
rect 38746 310536 38752 310548
rect 3384 310508 38752 310536
rect 3384 310496 3390 310508
rect 38746 310496 38752 310508
rect 38804 310496 38810 310548
rect 550266 307708 550272 307760
rect 550324 307748 550330 307760
rect 580166 307748 580172 307760
rect 550324 307720 580172 307748
rect 550324 307708 550330 307720
rect 580166 307708 580172 307720
rect 580224 307708 580230 307760
rect 16482 306280 16488 306332
rect 16540 306320 16546 306332
rect 38746 306320 38752 306332
rect 16540 306292 38752 306320
rect 16540 306280 16546 306292
rect 38746 306280 38752 306292
rect 38804 306280 38810 306332
rect 2774 304988 2780 305040
rect 2832 305028 2838 305040
rect 5350 305028 5356 305040
rect 2832 305000 5356 305028
rect 2832 304988 2838 305000
rect 5350 304988 5356 305000
rect 5408 304988 5414 305040
rect 556154 302336 556160 302388
rect 556212 302376 556218 302388
rect 559650 302376 559656 302388
rect 556212 302348 559656 302376
rect 556212 302336 556218 302348
rect 559650 302336 559656 302348
rect 559708 302336 559714 302388
rect 577498 302268 577504 302320
rect 577556 302308 577562 302320
rect 580810 302308 580816 302320
rect 577556 302280 580816 302308
rect 577556 302268 577562 302280
rect 580810 302268 580816 302280
rect 580868 302268 580874 302320
rect 550266 302200 550272 302252
rect 550324 302240 550330 302252
rect 580166 302240 580172 302252
rect 550324 302212 580172 302240
rect 550324 302200 550330 302212
rect 580166 302200 580172 302212
rect 580224 302200 580230 302252
rect 553118 299548 553124 299600
rect 553176 299588 553182 299600
rect 556154 299588 556160 299600
rect 553176 299560 556160 299588
rect 553176 299548 553182 299560
rect 556154 299548 556160 299560
rect 556212 299548 556218 299600
rect 550358 296692 550364 296744
rect 550416 296732 550422 296744
rect 579614 296732 579620 296744
rect 550416 296704 579620 296732
rect 550416 296692 550422 296704
rect 579614 296692 579620 296704
rect 579672 296692 579678 296744
rect 3326 295264 3332 295316
rect 3384 295304 3390 295316
rect 21450 295304 21456 295316
rect 3384 295276 21456 295304
rect 3384 295264 3390 295276
rect 21450 295264 21456 295276
rect 21508 295264 21514 295316
rect 35158 293904 35164 293956
rect 35216 293944 35222 293956
rect 38746 293944 38752 293956
rect 35216 293916 38752 293944
rect 35216 293904 35222 293916
rect 38746 293904 38752 293916
rect 38804 293904 38810 293956
rect 547690 292544 547696 292596
rect 547748 292584 547754 292596
rect 579798 292584 579804 292596
rect 547748 292556 579804 292584
rect 547748 292544 547754 292556
rect 579798 292544 579804 292556
rect 579856 292544 579862 292596
rect 3142 289824 3148 289876
rect 3200 289864 3206 289876
rect 11698 289864 11704 289876
rect 3200 289836 11704 289864
rect 3200 289824 3206 289836
rect 11698 289824 11704 289836
rect 11756 289824 11762 289876
rect 546218 287648 546224 287700
rect 546276 287688 546282 287700
rect 553118 287688 553124 287700
rect 546276 287660 553124 287688
rect 546276 287648 546282 287660
rect 553118 287648 553124 287660
rect 553176 287648 553182 287700
rect 563330 287648 563336 287700
rect 563388 287688 563394 287700
rect 577498 287688 577504 287700
rect 563388 287660 577504 287688
rect 563388 287648 563394 287660
rect 577498 287648 577504 287660
rect 577556 287648 577562 287700
rect 550542 287036 550548 287088
rect 550600 287076 550606 287088
rect 579614 287076 579620 287088
rect 550600 287048 579620 287076
rect 550600 287036 550606 287048
rect 579614 287036 579620 287048
rect 579672 287036 579678 287088
rect 561030 284316 561036 284368
rect 561088 284356 561094 284368
rect 563330 284356 563336 284368
rect 561088 284328 563336 284356
rect 561088 284316 561094 284328
rect 563330 284316 563336 284328
rect 563388 284316 563394 284368
rect 14458 284248 14464 284300
rect 14516 284288 14522 284300
rect 38746 284288 38752 284300
rect 14516 284260 38752 284288
rect 14516 284248 14522 284260
rect 38746 284248 38752 284260
rect 38804 284248 38810 284300
rect 547782 284248 547788 284300
rect 547840 284288 547846 284300
rect 579614 284288 579620 284300
rect 547840 284260 579620 284288
rect 547840 284248 547846 284260
rect 579614 284248 579620 284260
rect 579672 284248 579678 284300
rect 3326 280440 3332 280492
rect 3384 280480 3390 280492
rect 9490 280480 9496 280492
rect 3384 280452 9496 280480
rect 3384 280440 3390 280452
rect 9490 280440 9496 280452
rect 9548 280440 9554 280492
rect 37550 280100 37556 280152
rect 37608 280140 37614 280152
rect 39298 280140 39304 280152
rect 37608 280112 39304 280140
rect 37608 280100 37614 280112
rect 39298 280100 39304 280112
rect 39356 280100 39362 280152
rect 544930 278740 544936 278792
rect 544988 278780 544994 278792
rect 553302 278780 553308 278792
rect 544988 278752 553308 278780
rect 544988 278740 544994 278752
rect 553302 278740 553308 278752
rect 553360 278740 553366 278792
rect 553026 278672 553032 278724
rect 553084 278712 553090 278724
rect 579982 278712 579988 278724
rect 553084 278684 579988 278712
rect 553084 278672 553090 278684
rect 579982 278672 579988 278684
rect 580040 278672 580046 278724
rect 544746 275612 544752 275664
rect 544804 275652 544810 275664
rect 550450 275652 550456 275664
rect 544804 275624 550456 275652
rect 544804 275612 544810 275624
rect 550450 275612 550456 275624
rect 550508 275612 550514 275664
rect 39390 275340 39396 275392
rect 39448 275380 39454 275392
rect 40862 275380 40868 275392
rect 39448 275352 40868 275380
rect 39448 275340 39454 275352
rect 40862 275340 40868 275352
rect 40920 275340 40926 275392
rect 3326 274660 3332 274712
rect 3384 274700 3390 274712
rect 10870 274700 10876 274712
rect 3384 274672 10876 274700
rect 3384 274660 3390 274672
rect 10870 274660 10876 274672
rect 10928 274660 10934 274712
rect 553302 274592 553308 274644
rect 553360 274632 553366 274644
rect 580166 274632 580172 274644
rect 553360 274604 580172 274632
rect 553360 274592 553366 274604
rect 580166 274592 580172 274604
rect 580224 274592 580230 274644
rect 554774 273912 554780 273964
rect 554832 273952 554838 273964
rect 561030 273952 561036 273964
rect 554832 273924 561036 273952
rect 554832 273912 554838 273924
rect 561030 273912 561036 273924
rect 561088 273912 561094 273964
rect 553026 270716 553032 270768
rect 553084 270756 553090 270768
rect 554774 270756 554780 270768
rect 553084 270728 554780 270756
rect 553084 270716 553090 270728
rect 554774 270716 554780 270728
rect 554832 270716 554838 270768
rect 6546 270444 6552 270496
rect 6604 270484 6610 270496
rect 38746 270484 38752 270496
rect 6604 270456 38752 270484
rect 6604 270444 6610 270456
rect 38746 270444 38752 270456
rect 38804 270444 38810 270496
rect 546310 266976 546316 267028
rect 546368 267016 546374 267028
rect 553026 267016 553032 267028
rect 546368 266988 553032 267016
rect 546368 266976 546374 266988
rect 553026 266976 553032 266988
rect 553084 266976 553090 267028
rect 3142 266092 3148 266144
rect 3200 266132 3206 266144
rect 9582 266132 9588 266144
rect 3200 266104 9588 266132
rect 3200 266092 3206 266104
rect 9582 266092 9588 266104
rect 9640 266092 9646 266144
rect 546402 265684 546408 265736
rect 546460 265724 546466 265736
rect 556890 265724 556896 265736
rect 546460 265696 556896 265724
rect 546460 265684 546466 265696
rect 556890 265684 556896 265696
rect 556948 265684 556954 265736
rect 547046 265616 547052 265668
rect 547104 265656 547110 265668
rect 563054 265656 563060 265668
rect 547104 265628 563060 265656
rect 547104 265616 547110 265628
rect 563054 265616 563060 265628
rect 563112 265616 563118 265668
rect 3142 260176 3148 260228
rect 3200 260216 3206 260228
rect 9582 260216 9588 260228
rect 3200 260188 9588 260216
rect 3200 260176 3206 260188
rect 9582 260176 9588 260188
rect 9640 260176 9646 260228
rect 563054 260108 563060 260160
rect 563112 260148 563118 260160
rect 579798 260148 579804 260160
rect 563112 260120 579804 260148
rect 563112 260108 563118 260120
rect 579798 260108 579804 260120
rect 579856 260108 579862 260160
rect 551922 258068 551928 258120
rect 551980 258108 551986 258120
rect 580166 258108 580172 258120
rect 551980 258080 580172 258108
rect 551980 258068 551986 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 544746 255280 544752 255332
rect 544804 255320 544810 255332
rect 550450 255320 550456 255332
rect 544804 255292 550456 255320
rect 544804 255280 544810 255292
rect 550450 255280 550456 255292
rect 550508 255280 550514 255332
rect 556890 251812 556896 251864
rect 556948 251852 556954 251864
rect 572714 251852 572720 251864
rect 556948 251824 572720 251852
rect 556948 251812 556954 251824
rect 572714 251812 572720 251824
rect 572772 251812 572778 251864
rect 37550 251200 37556 251252
rect 37608 251240 37614 251252
rect 38746 251240 38752 251252
rect 37608 251212 38752 251240
rect 37608 251200 37614 251212
rect 38746 251200 38752 251212
rect 38804 251200 38810 251252
rect 572714 249704 572720 249756
rect 572772 249744 572778 249756
rect 579614 249744 579620 249756
rect 572772 249716 579620 249744
rect 572772 249704 572778 249716
rect 579614 249704 579620 249716
rect 579672 249704 579678 249756
rect 37642 248072 37648 248124
rect 37700 248112 37706 248124
rect 38838 248112 38844 248124
rect 37700 248084 38844 248112
rect 37700 248072 37706 248084
rect 38838 248072 38844 248084
rect 38896 248072 38902 248124
rect 544746 247052 544752 247104
rect 544804 247092 544810 247104
rect 553026 247092 553032 247104
rect 544804 247064 553032 247092
rect 544804 247052 544810 247064
rect 553026 247052 553032 247064
rect 553084 247052 553090 247104
rect 3602 246100 3608 246152
rect 3660 246140 3666 246152
rect 8110 246140 8116 246152
rect 3660 246112 8116 246140
rect 3660 246100 3666 246112
rect 8110 246100 8116 246112
rect 8168 246100 8174 246152
rect 11698 244196 11704 244248
rect 11756 244236 11762 244248
rect 38746 244236 38752 244248
rect 11756 244208 38752 244236
rect 11756 244196 11762 244208
rect 38746 244196 38752 244208
rect 38804 244196 38810 244248
rect 544746 242904 544752 242956
rect 544804 242944 544810 242956
rect 561030 242944 561036 242956
rect 544804 242916 561036 242944
rect 544804 242904 544810 242916
rect 561030 242904 561036 242916
rect 561088 242904 561094 242956
rect 3602 241068 3608 241120
rect 3660 241108 3666 241120
rect 9122 241108 9128 241120
rect 3660 241080 9128 241108
rect 3660 241068 3666 241080
rect 9122 241068 9128 241080
rect 9180 241068 9186 241120
rect 37734 240048 37740 240100
rect 37792 240088 37798 240100
rect 38746 240088 38752 240100
rect 37792 240060 38752 240088
rect 37792 240048 37798 240060
rect 38746 240048 38752 240060
rect 38804 240048 38810 240100
rect 545666 240048 545672 240100
rect 545724 240088 545730 240100
rect 580166 240088 580172 240100
rect 545724 240060 580172 240088
rect 545724 240048 545730 240060
rect 580166 240048 580172 240060
rect 580224 240048 580230 240100
rect 544746 237396 544752 237448
rect 544804 237436 544810 237448
rect 551186 237436 551192 237448
rect 544804 237408 551192 237436
rect 544804 237396 544810 237408
rect 551186 237396 551192 237408
rect 551244 237396 551250 237448
rect 3602 236172 3608 236224
rect 3660 236212 3666 236224
rect 7834 236212 7840 236224
rect 3660 236184 7840 236212
rect 3660 236172 3666 236184
rect 7834 236172 7840 236184
rect 7892 236172 7898 236224
rect 21358 234540 21364 234592
rect 21416 234580 21422 234592
rect 38746 234580 38752 234592
rect 21416 234552 38752 234580
rect 21416 234540 21422 234552
rect 38746 234540 38752 234552
rect 38804 234540 38810 234592
rect 553026 234540 553032 234592
rect 553084 234580 553090 234592
rect 579982 234580 579988 234592
rect 553084 234552 579988 234580
rect 553084 234540 553090 234552
rect 579982 234540 579988 234552
rect 580040 234540 580046 234592
rect 544470 229780 544476 229832
rect 544528 229820 544534 229832
rect 547414 229820 547420 229832
rect 544528 229792 547420 229820
rect 544528 229780 544534 229792
rect 547414 229780 547420 229792
rect 547472 229780 547478 229832
rect 574002 229100 574008 229152
rect 574060 229140 574066 229152
rect 580166 229140 580172 229152
rect 574060 229112 580172 229140
rect 574060 229100 574066 229112
rect 580166 229100 580172 229112
rect 580224 229100 580230 229152
rect 3142 226312 3148 226364
rect 3200 226352 3206 226364
rect 6546 226352 6552 226364
rect 3200 226324 6552 226352
rect 3200 226312 3206 226324
rect 6546 226312 6552 226324
rect 6604 226312 6610 226364
rect 544746 224952 544752 225004
rect 544804 224992 544810 225004
rect 553118 224992 553124 225004
rect 544804 224964 553124 224992
rect 544804 224952 544810 224964
rect 553118 224952 553124 224964
rect 553176 224952 553182 225004
rect 570598 223252 570604 223304
rect 570656 223292 570662 223304
rect 574002 223292 574008 223304
rect 570656 223264 574008 223292
rect 570656 223252 570662 223264
rect 574002 223252 574008 223264
rect 574060 223252 574066 223304
rect 3142 220804 3148 220856
rect 3200 220844 3206 220856
rect 38838 220844 38844 220856
rect 3200 220816 38844 220844
rect 3200 220804 3206 220816
rect 38838 220804 38844 220816
rect 38896 220804 38902 220856
rect 544746 219444 544752 219496
rect 544804 219484 544810 219496
rect 553026 219484 553032 219496
rect 544804 219456 553032 219484
rect 544804 219444 544810 219456
rect 553026 219444 553032 219456
rect 553084 219444 553090 219496
rect 560938 219376 560944 219428
rect 560996 219416 561002 219428
rect 579798 219416 579804 219428
rect 560996 219388 579804 219416
rect 560996 219376 561002 219388
rect 579798 219376 579804 219388
rect 579856 219376 579862 219428
rect 574738 215228 574744 215280
rect 574796 215268 574802 215280
rect 580166 215268 580172 215280
rect 574796 215240 580172 215268
rect 574796 215228 574802 215240
rect 580166 215228 580172 215240
rect 580224 215228 580230 215280
rect 3602 212440 3608 212492
rect 3660 212480 3666 212492
rect 33778 212480 33784 212492
rect 3660 212452 33784 212480
rect 3660 212440 3666 212452
rect 33778 212440 33784 212452
rect 33836 212440 33842 212492
rect 3050 211284 3056 211336
rect 3108 211324 3114 211336
rect 3602 211324 3608 211336
rect 3108 211296 3608 211324
rect 3108 211284 3114 211296
rect 3602 211284 3608 211296
rect 3660 211284 3666 211336
rect 544470 211148 544476 211200
rect 544528 211188 544534 211200
rect 547414 211188 547420 211200
rect 544528 211160 547420 211188
rect 544528 211148 544534 211160
rect 547414 211148 547420 211160
rect 547472 211148 547478 211200
rect 553118 209720 553124 209772
rect 553176 209760 553182 209772
rect 579982 209760 579988 209772
rect 553176 209732 579988 209760
rect 553176 209720 553182 209732
rect 579982 209720 579988 209732
rect 580040 209720 580046 209772
rect 553394 209040 553400 209092
rect 553452 209080 553458 209092
rect 570598 209080 570604 209092
rect 553452 209052 570604 209080
rect 553452 209040 553458 209052
rect 570598 209040 570604 209052
rect 570656 209040 570662 209092
rect 9214 208292 9220 208344
rect 9272 208332 9278 208344
rect 38838 208332 38844 208344
rect 9272 208304 38844 208332
rect 9272 208292 9278 208304
rect 38838 208292 38844 208304
rect 38896 208292 38902 208344
rect 544746 208292 544752 208344
rect 544804 208332 544810 208344
rect 564434 208332 564440 208344
rect 544804 208304 564440 208332
rect 544804 208292 544810 208304
rect 564434 208292 564440 208304
rect 564492 208292 564498 208344
rect 551094 205640 551100 205692
rect 551152 205680 551158 205692
rect 553394 205680 553400 205692
rect 551152 205652 553400 205680
rect 551152 205640 551158 205652
rect 553394 205640 553400 205652
rect 553452 205640 553458 205692
rect 3878 201424 3884 201476
rect 3936 201464 3942 201476
rect 5442 201464 5448 201476
rect 3936 201436 5448 201464
rect 3936 201424 3942 201436
rect 5442 201424 5448 201436
rect 5500 201424 5506 201476
rect 553026 200064 553032 200116
rect 553084 200104 553090 200116
rect 580166 200104 580172 200116
rect 553084 200076 580172 200104
rect 553084 200064 553090 200076
rect 580166 200064 580172 200076
rect 580224 200064 580230 200116
rect 3142 196664 3148 196716
rect 3200 196704 3206 196716
rect 9122 196704 9128 196716
rect 3200 196676 9128 196704
rect 3200 196664 3206 196676
rect 9122 196664 9128 196676
rect 9180 196664 9186 196716
rect 549070 195984 549076 196036
rect 549128 196024 549134 196036
rect 551094 196024 551100 196036
rect 549128 195996 551100 196024
rect 549128 195984 549134 195996
rect 551094 195984 551100 195996
rect 551152 195984 551158 196036
rect 5442 194488 5448 194540
rect 5500 194528 5506 194540
rect 8110 194528 8116 194540
rect 5500 194500 8116 194528
rect 5500 194488 5506 194500
rect 8110 194488 8116 194500
rect 8168 194488 8174 194540
rect 547414 194488 547420 194540
rect 547472 194528 547478 194540
rect 580166 194528 580172 194540
rect 547472 194500 580172 194528
rect 547472 194488 547478 194500
rect 580166 194488 580172 194500
rect 580224 194488 580230 194540
rect 11698 193196 11704 193248
rect 11756 193236 11762 193248
rect 38838 193236 38844 193248
rect 11756 193208 38844 193236
rect 11756 193196 11762 193208
rect 38838 193196 38844 193208
rect 38896 193196 38902 193248
rect 554130 190408 554136 190460
rect 554188 190448 554194 190460
rect 579614 190448 579620 190460
rect 554188 190420 579620 190448
rect 554188 190408 554194 190420
rect 579614 190408 579620 190420
rect 579672 190408 579678 190460
rect 37826 190068 37832 190120
rect 37884 190108 37890 190120
rect 39482 190108 39488 190120
rect 37884 190080 39488 190108
rect 37884 190068 37890 190080
rect 39482 190068 39488 190080
rect 39540 190068 39546 190120
rect 544470 189524 544476 189576
rect 544528 189564 544534 189576
rect 546402 189564 546408 189576
rect 544528 189536 546408 189564
rect 544528 189524 544534 189536
rect 546402 189524 546408 189536
rect 546460 189524 546466 189576
rect 3142 186600 3148 186652
rect 3200 186640 3206 186652
rect 7834 186640 7840 186652
rect 3200 186612 7840 186640
rect 3200 186600 3206 186612
rect 7834 186600 7840 186612
rect 7892 186600 7898 186652
rect 3050 184900 3056 184952
rect 3108 184940 3114 184952
rect 38838 184940 38844 184952
rect 3108 184912 38844 184940
rect 3108 184900 3114 184912
rect 38838 184900 38844 184912
rect 38896 184900 38902 184952
rect 546402 184900 546408 184952
rect 546460 184940 546466 184952
rect 546460 184912 547874 184940
rect 546460 184900 546466 184912
rect 547846 184872 547874 184912
rect 549806 184872 549812 184884
rect 547846 184844 549812 184872
rect 549806 184832 549812 184844
rect 549864 184832 549870 184884
rect 552842 184832 552848 184884
rect 552900 184872 552906 184884
rect 580166 184872 580172 184884
rect 552900 184844 580172 184872
rect 552900 184832 552906 184844
rect 580166 184832 580172 184844
rect 580224 184832 580230 184884
rect 544746 183540 544752 183592
rect 544804 183580 544810 183592
rect 565078 183580 565084 183592
rect 544804 183552 565084 183580
rect 544804 183540 544810 183552
rect 565078 183540 565084 183552
rect 565136 183540 565142 183592
rect 3142 182112 3148 182164
rect 3200 182152 3206 182164
rect 10686 182152 10692 182164
rect 3200 182124 10692 182152
rect 3200 182112 3206 182124
rect 10686 182112 10692 182124
rect 10744 182112 10750 182164
rect 546402 180820 546408 180872
rect 546460 180860 546466 180872
rect 549070 180860 549076 180872
rect 546460 180832 549076 180860
rect 546460 180820 546466 180832
rect 549070 180820 549076 180832
rect 549128 180820 549134 180872
rect 548610 180752 548616 180804
rect 548668 180792 548674 180804
rect 579982 180792 579988 180804
rect 548668 180764 579988 180792
rect 548668 180752 548674 180764
rect 579982 180752 579988 180764
rect 580040 180752 580046 180804
rect 543826 180548 543832 180600
rect 543884 180588 543890 180600
rect 546678 180588 546684 180600
rect 543884 180560 546684 180588
rect 543884 180548 543890 180560
rect 546678 180548 546684 180560
rect 546736 180548 546742 180600
rect 549806 178032 549812 178084
rect 549864 178072 549870 178084
rect 549864 178044 550680 178072
rect 549864 178032 549870 178044
rect 550652 178004 550680 178044
rect 554682 178004 554688 178016
rect 550652 177976 554688 178004
rect 554682 177964 554688 177976
rect 554740 177964 554746 178016
rect 3050 176944 3056 176996
rect 3108 176984 3114 176996
rect 6730 176984 6736 176996
rect 3108 176956 6736 176984
rect 3108 176944 3114 176956
rect 6730 176944 6736 176956
rect 6788 176944 6794 176996
rect 13078 176604 13084 176656
rect 13136 176644 13142 176656
rect 38838 176644 38844 176656
rect 13136 176616 38844 176644
rect 13136 176604 13142 176616
rect 38838 176604 38844 176616
rect 38896 176604 38902 176656
rect 544746 176604 544752 176656
rect 544804 176644 544810 176656
rect 559558 176644 559564 176656
rect 544804 176616 559564 176644
rect 544804 176604 544810 176616
rect 559558 176604 559564 176616
rect 559616 176604 559622 176656
rect 550450 175176 550456 175228
rect 550508 175216 550514 175228
rect 579614 175216 579620 175228
rect 550508 175188 579620 175216
rect 550508 175176 550514 175188
rect 579614 175176 579620 175188
rect 579672 175176 579678 175228
rect 8110 173816 8116 173868
rect 8168 173856 8174 173868
rect 12066 173856 12072 173868
rect 8168 173828 12072 173856
rect 8168 173816 8174 173828
rect 12066 173816 12072 173828
rect 12124 173816 12130 173868
rect 554774 172932 554780 172984
rect 554832 172972 554838 172984
rect 558914 172972 558920 172984
rect 554832 172944 558920 172972
rect 554832 172932 554838 172944
rect 558914 172932 558920 172944
rect 558972 172932 558978 172984
rect 3878 172456 3884 172508
rect 3936 172496 3942 172508
rect 5442 172496 5448 172508
rect 3936 172468 5448 172496
rect 3936 172456 3942 172468
rect 5442 172456 5448 172468
rect 5500 172456 5506 172508
rect 3050 172116 3056 172168
rect 3108 172156 3114 172168
rect 9214 172156 9220 172168
rect 3108 172128 9220 172156
rect 3108 172116 3114 172128
rect 9214 172116 9220 172128
rect 9272 172116 9278 172168
rect 545666 171776 545672 171828
rect 545724 171816 545730 171828
rect 580902 171816 580908 171828
rect 545724 171788 580908 171816
rect 545724 171776 545730 171788
rect 580902 171776 580908 171788
rect 580960 171776 580966 171828
rect 544470 171232 544476 171284
rect 544528 171272 544534 171284
rect 547414 171272 547420 171284
rect 544528 171244 547420 171272
rect 544528 171232 544534 171244
rect 547414 171232 547420 171244
rect 547472 171232 547478 171284
rect 558914 170348 558920 170400
rect 558972 170388 558978 170400
rect 569678 170388 569684 170400
rect 558972 170360 569684 170388
rect 558972 170348 558978 170360
rect 569678 170348 569684 170360
rect 569736 170348 569742 170400
rect 9582 168308 9588 168360
rect 9640 168348 9646 168360
rect 38838 168348 38844 168360
rect 9640 168320 38844 168348
rect 9640 168308 9646 168320
rect 38838 168308 38844 168320
rect 38896 168308 38902 168360
rect 543826 167220 543832 167272
rect 543884 167260 543890 167272
rect 546586 167260 546592 167272
rect 543884 167232 546592 167260
rect 543884 167220 543890 167232
rect 546586 167220 546592 167232
rect 546644 167220 546650 167272
rect 569678 167016 569684 167068
rect 569736 167056 569742 167068
rect 569736 167028 571380 167056
rect 569736 167016 569742 167028
rect 571352 166988 571380 167028
rect 574738 166988 574744 167000
rect 571352 166960 574744 166988
rect 574738 166948 574744 166960
rect 574796 166948 574802 167000
rect 12066 166540 12072 166592
rect 12124 166580 12130 166592
rect 14458 166580 14464 166592
rect 12124 166552 14464 166580
rect 12124 166540 12130 166552
rect 14458 166540 14464 166552
rect 14516 166540 14522 166592
rect 5442 165520 5448 165572
rect 5500 165560 5506 165572
rect 8110 165560 8116 165572
rect 5500 165532 8116 165560
rect 5500 165520 5506 165532
rect 8110 165520 8116 165532
rect 8168 165520 8174 165572
rect 547782 164228 547788 164280
rect 547840 164268 547846 164280
rect 579982 164268 579988 164280
rect 547840 164240 579988 164268
rect 547840 164228 547846 164240
rect 579982 164228 579988 164240
rect 580040 164228 580046 164280
rect 2774 162460 2780 162512
rect 2832 162500 2838 162512
rect 5074 162500 5080 162512
rect 2832 162472 5080 162500
rect 2832 162460 2838 162472
rect 5074 162460 5080 162472
rect 5132 162460 5138 162512
rect 17862 161440 17868 161492
rect 17920 161480 17926 161492
rect 38838 161480 38844 161492
rect 17920 161452 38844 161480
rect 17920 161440 17926 161452
rect 38838 161440 38844 161452
rect 38896 161440 38902 161492
rect 574738 160080 574744 160132
rect 574796 160120 574802 160132
rect 574796 160092 576854 160120
rect 574796 160080 574802 160092
rect 576826 160052 576854 160092
rect 580166 160052 580172 160064
rect 576826 160024 580172 160052
rect 580166 160012 580172 160024
rect 580224 160012 580230 160064
rect 544746 158652 544752 158704
rect 544804 158692 544810 158704
rect 556798 158692 556804 158704
rect 544804 158664 556804 158692
rect 544804 158652 544810 158664
rect 556798 158652 556804 158664
rect 556856 158652 556862 158704
rect 14458 155864 14464 155916
rect 14516 155904 14522 155916
rect 15194 155904 15200 155916
rect 14516 155876 15200 155904
rect 14516 155864 14522 155876
rect 15194 155864 15200 155876
rect 15252 155864 15258 155916
rect 565078 155864 565084 155916
rect 565136 155904 565142 155916
rect 579614 155904 579620 155916
rect 565136 155876 579620 155904
rect 565136 155864 565142 155876
rect 579614 155864 579620 155876
rect 579672 155864 579678 155916
rect 3786 153144 3792 153196
rect 3844 153184 3850 153196
rect 5350 153184 5356 153196
rect 3844 153156 5356 153184
rect 3844 153144 3850 153156
rect 5350 153144 5356 153156
rect 5408 153144 5414 153196
rect 15194 152056 15200 152108
rect 15252 152096 15258 152108
rect 17218 152096 17224 152108
rect 15252 152068 17224 152096
rect 15252 152056 15258 152068
rect 17218 152056 17224 152068
rect 17276 152056 17282 152108
rect 548610 149064 548616 149116
rect 548668 149104 548674 149116
rect 579614 149104 579620 149116
rect 548668 149076 579620 149104
rect 548668 149064 548674 149076
rect 579614 149064 579620 149076
rect 579672 149064 579678 149116
rect 3418 147568 3424 147620
rect 3476 147608 3482 147620
rect 25498 147608 25504 147620
rect 3476 147580 25504 147608
rect 3476 147568 3482 147580
rect 25498 147568 25504 147580
rect 25556 147568 25562 147620
rect 8110 144848 8116 144900
rect 8168 144888 8174 144900
rect 11790 144888 11796 144900
rect 8168 144860 11796 144888
rect 8168 144848 8174 144860
rect 11790 144848 11796 144860
rect 11848 144848 11854 144900
rect 17218 144848 17224 144900
rect 17276 144888 17282 144900
rect 18046 144888 18052 144900
rect 17276 144860 18052 144888
rect 17276 144848 17282 144860
rect 18046 144848 18052 144860
rect 18104 144848 18110 144900
rect 2774 142332 2780 142384
rect 2832 142372 2838 142384
rect 5074 142372 5080 142384
rect 2832 142344 5080 142372
rect 2832 142332 2838 142344
rect 5074 142332 5080 142344
rect 5132 142332 5138 142384
rect 18046 141108 18052 141160
rect 18104 141148 18110 141160
rect 21174 141148 21180 141160
rect 18104 141120 21180 141148
rect 18104 141108 18110 141120
rect 21174 141108 21180 141120
rect 21232 141108 21238 141160
rect 547322 140700 547328 140752
rect 547380 140740 547386 140752
rect 580166 140740 580172 140752
rect 547380 140712 580172 140740
rect 547380 140700 547386 140712
rect 580166 140700 580172 140712
rect 580224 140700 580230 140752
rect 5534 140292 5540 140344
rect 5592 140332 5598 140344
rect 8202 140332 8208 140344
rect 5592 140304 8208 140332
rect 5592 140292 5598 140304
rect 8202 140292 8208 140304
rect 8260 140292 8266 140344
rect 39942 139476 39948 139528
rect 40000 139516 40006 139528
rect 40954 139516 40960 139528
rect 40000 139488 40960 139516
rect 40000 139476 40006 139488
rect 40954 139476 40960 139488
rect 41012 139476 41018 139528
rect 3602 139408 3608 139460
rect 3660 139448 3666 139460
rect 3660 139420 4200 139448
rect 3660 139408 3666 139420
rect 4172 139380 4200 139420
rect 21174 139408 21180 139460
rect 21232 139448 21238 139460
rect 21232 139420 22140 139448
rect 21232 139408 21238 139420
rect 6086 139380 6092 139392
rect 4172 139352 6092 139380
rect 6086 139340 6092 139352
rect 6144 139340 6150 139392
rect 22112 139380 22140 139420
rect 24210 139380 24216 139392
rect 22112 139352 24216 139380
rect 24210 139340 24216 139352
rect 24268 139340 24274 139392
rect 8202 137844 8208 137896
rect 8260 137884 8266 137896
rect 9582 137884 9588 137896
rect 8260 137856 9588 137884
rect 8260 137844 8266 137856
rect 9582 137844 9588 137856
rect 9640 137844 9646 137896
rect 3418 137504 3424 137556
rect 3476 137544 3482 137556
rect 8110 137544 8116 137556
rect 3476 137516 8116 137544
rect 3476 137504 3482 137516
rect 8110 137504 8116 137516
rect 8168 137504 8174 137556
rect 11790 137504 11796 137556
rect 11848 137544 11854 137556
rect 14458 137544 14464 137556
rect 11848 137516 14464 137544
rect 11848 137504 11854 137516
rect 14458 137504 14464 137516
rect 14516 137504 14522 137556
rect 549070 135260 549076 135312
rect 549128 135300 549134 135312
rect 579614 135300 579620 135312
rect 549128 135272 579620 135300
rect 549128 135260 549134 135272
rect 579614 135260 579620 135272
rect 579672 135260 579678 135312
rect 33870 132404 33876 132456
rect 33928 132444 33934 132456
rect 38838 132444 38844 132456
rect 33928 132416 38844 132444
rect 33928 132404 33934 132416
rect 38838 132404 38844 132416
rect 38896 132404 38902 132456
rect 24210 131112 24216 131164
rect 24268 131152 24274 131164
rect 25498 131152 25504 131164
rect 24268 131124 25504 131152
rect 24268 131112 24274 131124
rect 25498 131112 25504 131124
rect 25556 131112 25562 131164
rect 6086 131044 6092 131096
rect 6144 131084 6150 131096
rect 8846 131084 8852 131096
rect 6144 131056 8852 131084
rect 6144 131044 6150 131056
rect 8846 131044 8852 131056
rect 8904 131044 8910 131096
rect 551186 131044 551192 131096
rect 551244 131084 551250 131096
rect 579798 131084 579804 131096
rect 551244 131056 579804 131084
rect 551244 131044 551250 131056
rect 579798 131044 579804 131056
rect 579856 131044 579862 131096
rect 3234 128256 3240 128308
rect 3292 128296 3298 128308
rect 10594 128296 10600 128308
rect 3292 128268 10600 128296
rect 3292 128256 3298 128268
rect 10594 128256 10600 128268
rect 10652 128256 10658 128308
rect 8846 126896 8852 126948
rect 8904 126936 8910 126948
rect 13078 126936 13084 126948
rect 8904 126908 13084 126936
rect 8904 126896 8910 126908
rect 13078 126896 13084 126908
rect 13136 126896 13142 126948
rect 14458 126896 14464 126948
rect 14516 126936 14522 126948
rect 15194 126936 15200 126948
rect 14516 126908 15200 126936
rect 14516 126896 14522 126908
rect 15194 126896 15200 126908
rect 15252 126896 15258 126948
rect 9582 126828 9588 126880
rect 9640 126868 9646 126880
rect 15838 126868 15844 126880
rect 9640 126840 15844 126868
rect 9640 126828 9646 126840
rect 15838 126828 15844 126840
rect 15896 126828 15902 126880
rect 3142 125604 3148 125656
rect 3200 125644 3206 125656
rect 3200 125616 4844 125644
rect 3200 125604 3206 125616
rect 3694 125536 3700 125588
rect 3752 125576 3758 125588
rect 4706 125576 4712 125588
rect 3752 125548 4712 125576
rect 3752 125536 3758 125548
rect 4706 125536 4712 125548
rect 4764 125536 4770 125588
rect 4816 125576 4844 125616
rect 5534 125576 5540 125588
rect 4816 125548 5540 125576
rect 5534 125536 5540 125548
rect 5592 125536 5598 125588
rect 15194 123156 15200 123208
rect 15252 123196 15258 123208
rect 17218 123196 17224 123208
rect 15252 123168 17224 123196
rect 15252 123156 15258 123168
rect 17218 123156 17224 123168
rect 17276 123156 17282 123208
rect 3602 122952 3608 123004
rect 3660 122992 3666 123004
rect 8202 122992 8208 123004
rect 3660 122964 8208 122992
rect 3660 122952 3666 122964
rect 8202 122952 8208 122964
rect 8260 122952 8266 123004
rect 13078 122204 13084 122256
rect 13136 122244 13142 122256
rect 14366 122244 14372 122256
rect 13136 122216 14372 122244
rect 13136 122204 13142 122216
rect 14366 122204 14372 122216
rect 14424 122204 14430 122256
rect 5534 120980 5540 121032
rect 5592 121020 5598 121032
rect 7466 121020 7472 121032
rect 5592 120992 7472 121020
rect 5592 120980 5598 120992
rect 7466 120980 7472 120992
rect 7524 120980 7530 121032
rect 552842 120096 552848 120148
rect 552900 120136 552906 120148
rect 580166 120136 580172 120148
rect 552900 120108 580172 120136
rect 552900 120096 552906 120108
rect 580166 120096 580172 120108
rect 580224 120096 580230 120148
rect 4706 118600 4712 118652
rect 4764 118640 4770 118652
rect 5534 118640 5540 118652
rect 4764 118612 5540 118640
rect 4764 118600 4770 118612
rect 5534 118600 5540 118612
rect 5592 118600 5598 118652
rect 3602 117308 3608 117360
rect 3660 117348 3666 117360
rect 12434 117348 12440 117360
rect 3660 117320 12440 117348
rect 3660 117308 3666 117320
rect 12434 117308 12440 117320
rect 12492 117308 12498 117360
rect 14366 117240 14372 117292
rect 14424 117280 14430 117292
rect 17310 117280 17316 117292
rect 14424 117252 17316 117280
rect 14424 117240 14430 117252
rect 17310 117240 17316 117252
rect 17368 117240 17374 117292
rect 561030 117240 561036 117292
rect 561088 117280 561094 117292
rect 579614 117280 579620 117292
rect 561088 117252 579620 117280
rect 561088 117240 561094 117252
rect 579614 117240 579620 117252
rect 579672 117240 579678 117292
rect 7466 117036 7472 117088
rect 7524 117076 7530 117088
rect 9582 117076 9588 117088
rect 7524 117048 9588 117076
rect 7524 117036 7530 117048
rect 9582 117036 9588 117048
rect 9640 117036 9646 117088
rect 12434 115744 12440 115796
rect 12492 115784 12498 115796
rect 16206 115784 16212 115796
rect 12492 115756 16212 115784
rect 12492 115744 12498 115756
rect 16206 115744 16212 115756
rect 16264 115744 16270 115796
rect 5534 115608 5540 115660
rect 5592 115648 5598 115660
rect 7466 115648 7472 115660
rect 5592 115620 7472 115648
rect 5592 115608 5598 115620
rect 7466 115608 7472 115620
rect 7524 115608 7530 115660
rect 25498 115132 25504 115184
rect 25556 115172 25562 115184
rect 27614 115172 27620 115184
rect 25556 115144 27620 115172
rect 25556 115132 25562 115144
rect 27614 115132 27620 115144
rect 27672 115132 27678 115184
rect 20622 114452 20628 114504
rect 20680 114492 20686 114504
rect 38838 114492 38844 114504
rect 20680 114464 38844 114492
rect 20680 114452 20686 114464
rect 38838 114452 38844 114464
rect 38896 114452 38902 114504
rect 544654 114452 544660 114504
rect 544712 114492 544718 114504
rect 558178 114492 558184 114504
rect 544712 114464 558184 114492
rect 544712 114452 544718 114464
rect 558178 114452 558184 114464
rect 558236 114452 558242 114504
rect 3050 113160 3056 113212
rect 3108 113200 3114 113212
rect 6086 113200 6092 113212
rect 3108 113172 6092 113200
rect 3108 113160 3114 113172
rect 6086 113160 6092 113172
rect 6144 113160 6150 113212
rect 9582 110440 9588 110492
rect 9640 110480 9646 110492
rect 9640 110452 11100 110480
rect 9640 110440 9646 110452
rect 11072 110412 11100 110452
rect 17310 110440 17316 110492
rect 17368 110480 17374 110492
rect 17368 110452 18000 110480
rect 17368 110440 17374 110452
rect 12434 110412 12440 110424
rect 11072 110384 12440 110412
rect 12434 110372 12440 110384
rect 12492 110372 12498 110424
rect 17972 110412 18000 110452
rect 27614 110440 27620 110492
rect 27672 110480 27678 110492
rect 29638 110480 29644 110492
rect 27672 110452 29644 110480
rect 27672 110440 27678 110452
rect 29638 110440 29644 110452
rect 29696 110440 29702 110492
rect 567746 110440 567752 110492
rect 567804 110480 567810 110492
rect 580166 110480 580172 110492
rect 567804 110452 580172 110480
rect 567804 110440 567810 110452
rect 580166 110440 580172 110452
rect 580224 110440 580230 110492
rect 20162 110412 20168 110424
rect 17972 110384 20168 110412
rect 20162 110372 20168 110384
rect 20220 110372 20226 110424
rect 7466 109624 7472 109676
rect 7524 109664 7530 109676
rect 10594 109664 10600 109676
rect 7524 109636 10600 109664
rect 7524 109624 7530 109636
rect 10594 109624 10600 109636
rect 10652 109624 10658 109676
rect 3326 109556 3332 109608
rect 3384 109596 3390 109608
rect 5350 109596 5356 109608
rect 3384 109568 5356 109596
rect 3384 109556 3390 109568
rect 5350 109556 5356 109568
rect 5408 109556 5414 109608
rect 10778 108944 10784 108996
rect 10836 108984 10842 108996
rect 38838 108984 38844 108996
rect 10836 108956 38844 108984
rect 10836 108944 10842 108956
rect 38838 108944 38844 108956
rect 38896 108944 38902 108996
rect 3142 108672 3148 108724
rect 3200 108712 3206 108724
rect 6638 108712 6644 108724
rect 3200 108684 6644 108712
rect 3200 108672 3206 108684
rect 6638 108672 6644 108684
rect 6696 108672 6702 108724
rect 16206 108264 16212 108316
rect 16264 108304 16270 108316
rect 19978 108304 19984 108316
rect 16264 108276 19984 108304
rect 16264 108264 16270 108276
rect 19978 108264 19984 108276
rect 20036 108264 20042 108316
rect 5350 107584 5356 107636
rect 5408 107624 5414 107636
rect 6638 107624 6644 107636
rect 5408 107596 6644 107624
rect 5408 107584 5414 107596
rect 6638 107584 6644 107596
rect 6696 107584 6702 107636
rect 12434 107584 12440 107636
rect 12492 107624 12498 107636
rect 17402 107624 17408 107636
rect 12492 107596 17408 107624
rect 12492 107584 12498 107596
rect 17402 107584 17408 107596
rect 17460 107584 17466 107636
rect 20162 107584 20168 107636
rect 20220 107624 20226 107636
rect 22830 107624 22836 107636
rect 20220 107596 22836 107624
rect 20220 107584 20226 107596
rect 22830 107584 22836 107596
rect 22888 107584 22894 107636
rect 17218 107516 17224 107568
rect 17276 107556 17282 107568
rect 20070 107556 20076 107568
rect 17276 107528 20076 107556
rect 17276 107516 17282 107528
rect 20070 107516 20076 107528
rect 20128 107516 20134 107568
rect 17402 104796 17408 104848
rect 17460 104836 17466 104848
rect 18322 104836 18328 104848
rect 17460 104808 18328 104836
rect 17460 104796 17466 104808
rect 18322 104796 18328 104808
rect 18380 104796 18386 104848
rect 543550 104116 543556 104168
rect 543608 104156 543614 104168
rect 567746 104156 567752 104168
rect 543608 104128 567752 104156
rect 543608 104116 543614 104128
rect 567746 104116 567752 104128
rect 567804 104116 567810 104168
rect 3326 103436 3332 103488
rect 3384 103476 3390 103488
rect 24118 103476 24124 103488
rect 3384 103448 24124 103476
rect 3384 103436 3390 103448
rect 24118 103436 24124 103448
rect 24176 103436 24182 103488
rect 6638 102620 6644 102672
rect 6696 102660 6702 102672
rect 7466 102660 7472 102672
rect 6696 102632 7472 102660
rect 6696 102620 6702 102632
rect 7466 102620 7472 102632
rect 7524 102620 7530 102672
rect 20070 102484 20076 102536
rect 20128 102524 20134 102536
rect 21542 102524 21548 102536
rect 20128 102496 21548 102524
rect 20128 102484 20134 102496
rect 21542 102484 21548 102496
rect 21600 102484 21606 102536
rect 578234 102144 578240 102196
rect 578292 102184 578298 102196
rect 580166 102184 580172 102196
rect 578292 102156 580172 102184
rect 578292 102144 578298 102156
rect 580166 102144 580172 102156
rect 580224 102144 580230 102196
rect 549990 102076 549996 102128
rect 550048 102116 550054 102128
rect 579614 102116 579620 102128
rect 550048 102088 579620 102116
rect 550048 102076 550054 102088
rect 579614 102076 579620 102088
rect 579672 102076 579678 102128
rect 18322 100988 18328 101040
rect 18380 101028 18386 101040
rect 21358 101028 21364 101040
rect 18380 101000 21364 101028
rect 18380 100988 18386 101000
rect 21358 100988 21364 101000
rect 21416 100988 21422 101040
rect 19978 100716 19984 100768
rect 20036 100756 20042 100768
rect 21450 100756 21456 100768
rect 20036 100728 21456 100756
rect 20036 100716 20042 100728
rect 21450 100716 21456 100728
rect 21508 100716 21514 100768
rect 21542 100580 21548 100632
rect 21600 100620 21606 100632
rect 22738 100620 22744 100632
rect 21600 100592 22744 100620
rect 21600 100580 21606 100592
rect 22738 100580 22744 100592
rect 22796 100580 22802 100632
rect 15838 99968 15844 100020
rect 15896 100008 15902 100020
rect 20714 100008 20720 100020
rect 15896 99980 20720 100008
rect 15896 99968 15902 99980
rect 20714 99968 20720 99980
rect 20772 99968 20778 100020
rect 22830 99084 22836 99136
rect 22888 99124 22894 99136
rect 24118 99124 24124 99136
rect 22888 99096 24124 99124
rect 22888 99084 22894 99096
rect 24118 99084 24124 99096
rect 24176 99084 24182 99136
rect 7466 99016 7472 99068
rect 7524 99056 7530 99068
rect 8846 99056 8852 99068
rect 7524 99028 8852 99056
rect 7524 99016 7530 99028
rect 8846 99016 8852 99028
rect 8904 99016 8910 99068
rect 10594 98812 10600 98864
rect 10652 98852 10658 98864
rect 11790 98852 11796 98864
rect 10652 98824 11796 98852
rect 10652 98812 10658 98824
rect 11790 98812 11796 98824
rect 11848 98812 11854 98864
rect 39114 97928 39120 97980
rect 39172 97968 39178 97980
rect 41138 97968 41144 97980
rect 39172 97940 41144 97968
rect 39172 97928 39178 97940
rect 41138 97928 41144 97940
rect 41196 97928 41202 97980
rect 566458 97248 566464 97300
rect 566516 97288 566522 97300
rect 578142 97288 578148 97300
rect 566516 97260 578148 97288
rect 566516 97248 566522 97260
rect 578142 97248 578148 97260
rect 578200 97248 578206 97300
rect 8846 96568 8852 96620
rect 8904 96608 8910 96620
rect 16482 96608 16488 96620
rect 8904 96580 16488 96608
rect 8904 96568 8910 96580
rect 16482 96568 16488 96580
rect 16540 96568 16546 96620
rect 20714 95140 20720 95192
rect 20772 95180 20778 95192
rect 22830 95180 22836 95192
rect 20772 95152 22836 95180
rect 20772 95140 20778 95152
rect 22830 95140 22836 95152
rect 22888 95140 22894 95192
rect 543366 95140 543372 95192
rect 543424 95180 543430 95192
rect 543734 95180 543740 95192
rect 543424 95152 543740 95180
rect 543424 95140 543430 95152
rect 543734 95140 543740 95152
rect 543792 95140 543798 95192
rect 563790 94460 563796 94512
rect 563848 94500 563854 94512
rect 580718 94500 580724 94512
rect 563848 94472 580724 94500
rect 563848 94460 563854 94472
rect 580718 94460 580724 94472
rect 580776 94460 580782 94512
rect 40954 93508 40960 93560
rect 41012 93548 41018 93560
rect 41598 93548 41604 93560
rect 41012 93520 41604 93548
rect 41012 93508 41018 93520
rect 41598 93508 41604 93520
rect 41656 93508 41662 93560
rect 2774 92760 2780 92812
rect 2832 92800 2838 92812
rect 5350 92800 5356 92812
rect 2832 92772 5356 92800
rect 2832 92760 2838 92772
rect 5350 92760 5356 92772
rect 5408 92760 5414 92812
rect 16574 92488 16580 92540
rect 16632 92528 16638 92540
rect 16632 92500 20760 92528
rect 16632 92488 16638 92500
rect 20732 92460 20760 92500
rect 25682 92460 25688 92472
rect 20732 92432 25688 92460
rect 25682 92420 25688 92432
rect 25740 92420 25746 92472
rect 38930 92012 38936 92064
rect 38988 92052 38994 92064
rect 41046 92052 41052 92064
rect 38988 92024 41052 92052
rect 38988 92012 38994 92024
rect 41046 92012 41052 92024
rect 41104 92012 41110 92064
rect 11790 91876 11796 91928
rect 11848 91916 11854 91928
rect 13722 91916 13728 91928
rect 11848 91888 13728 91916
rect 11848 91876 11854 91888
rect 13722 91876 13728 91888
rect 13780 91876 13786 91928
rect 22738 91060 22744 91112
rect 22796 91100 22802 91112
rect 22796 91072 23520 91100
rect 22796 91060 22802 91072
rect 23492 91032 23520 91072
rect 25498 91032 25504 91044
rect 23492 91004 25504 91032
rect 25498 90992 25504 91004
rect 25556 90992 25562 91044
rect 561766 89700 561772 89752
rect 561824 89740 561830 89752
rect 566458 89740 566464 89752
rect 561824 89712 566464 89740
rect 561824 89700 561830 89712
rect 566458 89700 566464 89712
rect 566516 89700 566522 89752
rect 13722 88340 13728 88392
rect 13780 88380 13786 88392
rect 13780 88352 13860 88380
rect 13780 88340 13786 88352
rect 13832 88312 13860 88352
rect 15194 88312 15200 88324
rect 13832 88284 15200 88312
rect 15194 88272 15200 88284
rect 15252 88272 15258 88324
rect 24118 88272 24124 88324
rect 24176 88312 24182 88324
rect 25590 88312 25596 88324
rect 24176 88284 25596 88312
rect 24176 88272 24182 88284
rect 25590 88272 25596 88284
rect 25648 88272 25654 88324
rect 29638 88272 29644 88324
rect 29696 88312 29702 88324
rect 32398 88312 32404 88324
rect 29696 88284 32404 88312
rect 29696 88272 29702 88284
rect 32398 88272 32404 88284
rect 32456 88272 32462 88324
rect 22830 86912 22836 86964
rect 22888 86952 22894 86964
rect 24118 86952 24124 86964
rect 22888 86924 24124 86952
rect 22888 86912 22894 86924
rect 24118 86912 24124 86924
rect 24176 86912 24182 86964
rect 544838 86232 544844 86284
rect 544896 86272 544902 86284
rect 563790 86272 563796 86284
rect 544896 86244 563796 86272
rect 544896 86232 544902 86244
rect 563790 86232 563796 86244
rect 563848 86232 563854 86284
rect 15194 85552 15200 85604
rect 15252 85592 15258 85604
rect 15252 85564 16574 85592
rect 15252 85552 15258 85564
rect 16546 85524 16574 85564
rect 558822 85552 558828 85604
rect 558880 85592 558886 85604
rect 561766 85592 561772 85604
rect 558880 85564 561772 85592
rect 558880 85552 558886 85564
rect 561766 85552 561772 85564
rect 561824 85552 561830 85604
rect 18598 85524 18604 85536
rect 16546 85496 18604 85524
rect 18598 85484 18604 85496
rect 18656 85484 18662 85536
rect 21450 84192 21456 84244
rect 21508 84232 21514 84244
rect 21508 84204 22140 84232
rect 21508 84192 21514 84204
rect 22112 84164 22140 84204
rect 551186 84192 551192 84244
rect 551244 84232 551250 84244
rect 558822 84232 558828 84244
rect 551244 84204 558828 84232
rect 551244 84192 551250 84204
rect 558822 84192 558828 84204
rect 558880 84192 558886 84244
rect 23934 84164 23940 84176
rect 22112 84136 23940 84164
rect 23934 84124 23940 84136
rect 23992 84124 23998 84176
rect 25682 83104 25688 83156
rect 25740 83144 25746 83156
rect 27522 83144 27528 83156
rect 25740 83116 27528 83144
rect 25740 83104 25746 83116
rect 27522 83104 27528 83116
rect 27580 83104 27586 83156
rect 3326 82832 3332 82884
rect 3384 82872 3390 82884
rect 3384 82844 21404 82872
rect 3384 82832 3390 82844
rect 21376 82804 21404 82844
rect 24854 82804 24860 82816
rect 21376 82776 24860 82804
rect 24854 82764 24860 82776
rect 24912 82764 24918 82816
rect 39850 82628 39856 82680
rect 39908 82668 39914 82680
rect 41322 82668 41328 82680
rect 39908 82640 41328 82668
rect 39908 82628 39914 82640
rect 41322 82628 41328 82640
rect 41380 82628 41386 82680
rect 40034 82356 40040 82408
rect 40092 82396 40098 82408
rect 41506 82396 41512 82408
rect 40092 82368 41512 82396
rect 40092 82356 40098 82368
rect 41506 82356 41512 82368
rect 41564 82356 41570 82408
rect 543826 81404 543832 81456
rect 543884 81444 543890 81456
rect 558178 81444 558184 81456
rect 543884 81416 558184 81444
rect 543884 81404 543890 81416
rect 558178 81404 558184 81416
rect 558236 81404 558242 81456
rect 545758 81336 545764 81388
rect 545816 81376 545822 81388
rect 580166 81376 580172 81388
rect 545816 81348 580172 81376
rect 545816 81336 545822 81348
rect 580166 81336 580172 81348
rect 580224 81336 580230 81388
rect 549530 79772 549536 79824
rect 549588 79812 549594 79824
rect 551186 79812 551192 79824
rect 549588 79784 551192 79812
rect 549588 79772 549594 79784
rect 551186 79772 551192 79784
rect 551244 79772 551250 79824
rect 23934 79364 23940 79416
rect 23992 79404 23998 79416
rect 25774 79404 25780 79416
rect 23992 79376 25780 79404
rect 23992 79364 23998 79376
rect 25774 79364 25780 79376
rect 25832 79364 25838 79416
rect 27522 79024 27528 79076
rect 27580 79064 27586 79076
rect 28994 79064 29000 79076
rect 27580 79036 29000 79064
rect 27580 79024 27586 79036
rect 28994 79024 29000 79036
rect 29052 79024 29058 79076
rect 2774 78684 2780 78736
rect 2832 78724 2838 78736
rect 5442 78724 5448 78736
rect 2832 78696 5448 78724
rect 2832 78684 2838 78696
rect 5442 78684 5448 78696
rect 5500 78684 5506 78736
rect 24854 78616 24860 78668
rect 24912 78656 24918 78668
rect 27246 78656 27252 78668
rect 24912 78628 27252 78656
rect 24912 78616 24918 78628
rect 27246 78616 27252 78628
rect 27304 78616 27310 78668
rect 32398 78616 32404 78668
rect 32456 78656 32462 78668
rect 36538 78656 36544 78668
rect 32456 78628 36544 78656
rect 32456 78616 32462 78628
rect 36538 78616 36544 78628
rect 36596 78616 36602 78668
rect 21358 77256 21364 77308
rect 21416 77296 21422 77308
rect 21416 77268 22140 77296
rect 21416 77256 21422 77268
rect 18598 77188 18604 77240
rect 18656 77228 18662 77240
rect 20622 77228 20628 77240
rect 18656 77200 20628 77228
rect 18656 77188 18662 77200
rect 20622 77188 20628 77200
rect 20680 77188 20686 77240
rect 22112 77228 22140 77268
rect 28994 77256 29000 77308
rect 29052 77296 29058 77308
rect 29052 77268 30420 77296
rect 29052 77256 29058 77268
rect 25406 77228 25412 77240
rect 22112 77200 25412 77228
rect 25406 77188 25412 77200
rect 25464 77188 25470 77240
rect 30392 77228 30420 77268
rect 33778 77228 33784 77240
rect 30392 77200 33784 77228
rect 33778 77188 33784 77200
rect 33836 77188 33842 77240
rect 25498 77052 25504 77104
rect 25556 77092 25562 77104
rect 26970 77092 26976 77104
rect 25556 77064 26976 77092
rect 25556 77052 25562 77064
rect 26970 77052 26976 77064
rect 27028 77052 27034 77104
rect 25590 75896 25596 75948
rect 25648 75936 25654 75948
rect 26878 75936 26884 75948
rect 25648 75908 26884 75936
rect 25648 75896 25654 75908
rect 26878 75896 26884 75908
rect 26936 75896 26942 75948
rect 549530 75936 549536 75948
rect 543752 75908 549536 75936
rect 27246 75828 27252 75880
rect 27304 75868 27310 75880
rect 30282 75868 30288 75880
rect 27304 75840 30288 75868
rect 27304 75828 27310 75840
rect 30282 75828 30288 75840
rect 30340 75828 30346 75880
rect 543642 75828 543648 75880
rect 543700 75868 543706 75880
rect 543752 75868 543780 75908
rect 549530 75896 549536 75908
rect 549588 75896 549594 75948
rect 543700 75840 543780 75868
rect 543700 75828 543706 75840
rect 24118 74536 24124 74588
rect 24176 74576 24182 74588
rect 24176 74548 24900 74576
rect 24176 74536 24182 74548
rect 3326 74468 3332 74520
rect 3384 74508 3390 74520
rect 10410 74508 10416 74520
rect 3384 74480 10416 74508
rect 3384 74468 3390 74480
rect 10410 74468 10416 74480
rect 10468 74468 10474 74520
rect 24872 74508 24900 74548
rect 27522 74508 27528 74520
rect 24872 74480 27528 74508
rect 27522 74468 27528 74480
rect 27580 74468 27586 74520
rect 39942 73652 39948 73704
rect 40000 73692 40006 73704
rect 41690 73692 41696 73704
rect 40000 73664 41696 73692
rect 40000 73652 40006 73664
rect 41690 73652 41696 73664
rect 41748 73652 41754 73704
rect 542262 73176 542268 73228
rect 542320 73216 542326 73228
rect 543550 73216 543556 73228
rect 542320 73188 543556 73216
rect 542320 73176 542326 73188
rect 543550 73176 543556 73188
rect 543608 73176 543614 73228
rect 25774 73108 25780 73160
rect 25832 73148 25838 73160
rect 27246 73148 27252 73160
rect 25832 73120 27252 73148
rect 25832 73108 25838 73120
rect 27246 73108 27252 73120
rect 27304 73108 27310 73160
rect 27522 71748 27528 71800
rect 27580 71788 27586 71800
rect 27580 71760 27660 71788
rect 27580 71748 27586 71760
rect 27632 71720 27660 71760
rect 29086 71720 29092 71732
rect 27632 71692 29092 71720
rect 29086 71680 29092 71692
rect 29144 71680 29150 71732
rect 27246 70456 27252 70508
rect 27304 70496 27310 70508
rect 31018 70496 31024 70508
rect 27304 70468 31024 70496
rect 27304 70456 27310 70468
rect 31018 70456 31024 70468
rect 31076 70456 31082 70508
rect 30374 69844 30380 69896
rect 30432 69884 30438 69896
rect 35158 69884 35164 69896
rect 30432 69856 35164 69884
rect 30432 69844 30438 69856
rect 35158 69844 35164 69856
rect 35216 69844 35222 69896
rect 25406 69028 25412 69080
rect 25464 69068 25470 69080
rect 25464 69040 26234 69068
rect 25464 69028 25470 69040
rect 26206 69000 26234 69040
rect 29086 69028 29092 69080
rect 29144 69068 29150 69080
rect 29144 69040 30420 69068
rect 29144 69028 29150 69040
rect 27614 69000 27620 69012
rect 26206 68972 27620 69000
rect 27614 68960 27620 68972
rect 27672 68960 27678 69012
rect 30392 69000 30420 69040
rect 32490 69000 32496 69012
rect 30392 68972 32496 69000
rect 32490 68960 32496 68972
rect 32548 68960 32554 69012
rect 543826 68960 543832 69012
rect 543884 69000 543890 69012
rect 554038 69000 554044 69012
rect 543884 68972 554044 69000
rect 543884 68960 543890 68972
rect 554038 68960 554044 68972
rect 554096 68960 554102 69012
rect 3326 68892 3332 68944
rect 3384 68932 3390 68944
rect 8018 68932 8024 68944
rect 3384 68904 8024 68932
rect 3384 68892 3390 68904
rect 8018 68892 8024 68904
rect 8076 68892 8082 68944
rect 20714 68280 20720 68332
rect 20772 68320 20778 68332
rect 29638 68320 29644 68332
rect 20772 68292 29644 68320
rect 20772 68280 20778 68292
rect 29638 68280 29644 68292
rect 29696 68280 29702 68332
rect 27614 67532 27620 67584
rect 27672 67572 27678 67584
rect 30282 67572 30288 67584
rect 27672 67544 30288 67572
rect 27672 67532 27678 67544
rect 30282 67532 30288 67544
rect 30340 67532 30346 67584
rect 575474 66240 575480 66292
rect 575532 66280 575538 66292
rect 578970 66280 578976 66292
rect 575532 66252 578976 66280
rect 575532 66240 575538 66252
rect 578970 66240 578976 66252
rect 579028 66240 579034 66292
rect 38838 64744 38844 64796
rect 38896 64784 38902 64796
rect 40954 64784 40960 64796
rect 38896 64756 40960 64784
rect 38896 64744 38902 64756
rect 40954 64744 40960 64756
rect 41012 64744 41018 64796
rect 31018 64132 31024 64184
rect 31076 64172 31082 64184
rect 32398 64172 32404 64184
rect 31076 64144 32404 64172
rect 31076 64132 31082 64144
rect 32398 64132 32404 64144
rect 32456 64132 32462 64184
rect 543826 64132 543832 64184
rect 543884 64172 543890 64184
rect 545942 64172 545948 64184
rect 543884 64144 545948 64172
rect 543884 64132 543890 64144
rect 545942 64132 545948 64144
rect 546000 64132 546006 64184
rect 2774 63996 2780 64048
rect 2832 64036 2838 64048
rect 4798 64036 4804 64048
rect 2832 64008 4804 64036
rect 2832 63996 2838 64008
rect 4798 63996 4804 64008
rect 4856 63996 4862 64048
rect 26970 63724 26976 63776
rect 27028 63764 27034 63776
rect 31478 63764 31484 63776
rect 27028 63736 31484 63764
rect 27028 63724 27034 63736
rect 31478 63724 31484 63736
rect 31536 63724 31542 63776
rect 35158 63520 35164 63572
rect 35216 63560 35222 63572
rect 35216 63532 35894 63560
rect 35216 63520 35222 63532
rect 35866 63492 35894 63532
rect 38102 63492 38108 63504
rect 35866 63464 38108 63492
rect 38102 63452 38108 63464
rect 38160 63452 38166 63504
rect 30282 62636 30288 62688
rect 30340 62676 30346 62688
rect 32306 62676 32312 62688
rect 30340 62648 32312 62676
rect 30340 62636 30346 62648
rect 32306 62636 32312 62648
rect 32364 62636 32370 62688
rect 575382 62132 575388 62144
rect 572732 62104 575388 62132
rect 571702 62024 571708 62076
rect 571760 62064 571766 62076
rect 572732 62064 572760 62104
rect 575382 62092 575388 62104
rect 575440 62092 575446 62144
rect 571760 62036 572760 62064
rect 571760 62024 571766 62036
rect 33778 60596 33784 60648
rect 33836 60636 33842 60648
rect 34514 60636 34520 60648
rect 33836 60608 34520 60636
rect 33836 60596 33842 60608
rect 34514 60596 34520 60608
rect 34572 60596 34578 60648
rect 26878 60188 26884 60240
rect 26936 60228 26942 60240
rect 31662 60228 31668 60240
rect 26936 60200 31668 60228
rect 26936 60188 26942 60200
rect 31662 60188 31668 60200
rect 31720 60188 31726 60240
rect 543826 59508 543832 59560
rect 543884 59548 543890 59560
rect 546494 59548 546500 59560
rect 543884 59520 546500 59548
rect 543884 59508 543890 59520
rect 546494 59508 546500 59520
rect 546552 59508 546558 59560
rect 3694 59372 3700 59424
rect 3752 59412 3758 59424
rect 38838 59412 38844 59424
rect 3752 59384 38844 59412
rect 3752 59372 3758 59384
rect 38838 59372 38844 59384
rect 38896 59372 38902 59424
rect 31478 59304 31484 59356
rect 31536 59344 31542 59356
rect 33134 59344 33140 59356
rect 31536 59316 33140 59344
rect 31536 59304 31542 59316
rect 33134 59304 33140 59316
rect 33192 59304 33198 59356
rect 567930 59304 567936 59356
rect 567988 59344 567994 59356
rect 571702 59344 571708 59356
rect 567988 59316 571708 59344
rect 567988 59304 567994 59316
rect 571702 59304 571708 59316
rect 571760 59304 571766 59356
rect 32306 57876 32312 57928
rect 32364 57916 32370 57928
rect 34422 57916 34428 57928
rect 32364 57888 34428 57916
rect 32364 57876 32370 57888
rect 34422 57876 34428 57888
rect 34480 57876 34486 57928
rect 31754 56584 31760 56636
rect 31812 56624 31818 56636
rect 31812 56596 33180 56624
rect 31812 56584 31818 56596
rect 33152 56556 33180 56596
rect 35618 56556 35624 56568
rect 33152 56528 35624 56556
rect 35618 56516 35624 56528
rect 35676 56516 35682 56568
rect 39206 56516 39212 56568
rect 39264 56556 39270 56568
rect 41230 56556 41236 56568
rect 39264 56528 41236 56556
rect 39264 56516 39270 56528
rect 41230 56516 41236 56528
rect 41288 56516 41294 56568
rect 33134 56108 33140 56160
rect 33192 56148 33198 56160
rect 36630 56148 36636 56160
rect 33192 56120 36636 56148
rect 33192 56108 33198 56120
rect 36630 56108 36636 56120
rect 36688 56108 36694 56160
rect 34514 55700 34520 55752
rect 34572 55740 34578 55752
rect 36814 55740 36820 55752
rect 34572 55712 36820 55740
rect 34572 55700 34578 55712
rect 36814 55700 36820 55712
rect 36872 55700 36878 55752
rect 541897 53839 541955 53845
rect 541897 53805 541909 53839
rect 541943 53836 541955 53839
rect 543826 53836 543832 53848
rect 541943 53808 543832 53836
rect 541943 53805 541955 53808
rect 541897 53799 541955 53805
rect 543826 53796 543832 53808
rect 543884 53796 543890 53848
rect 35618 53048 35624 53100
rect 35676 53088 35682 53100
rect 41414 53088 41420 53100
rect 35676 53060 41420 53088
rect 35676 53048 35682 53060
rect 41414 53048 41420 53060
rect 41472 53048 41478 53100
rect 564434 52776 564440 52828
rect 564492 52816 564498 52828
rect 567930 52816 567936 52828
rect 564492 52788 567936 52816
rect 564492 52776 564498 52788
rect 567930 52776 567936 52788
rect 567988 52776 567994 52828
rect 38102 52436 38108 52488
rect 38160 52476 38166 52488
rect 39206 52476 39212 52488
rect 38160 52448 39212 52476
rect 38160 52436 38166 52448
rect 39206 52436 39212 52448
rect 39264 52436 39270 52488
rect 567838 52368 567844 52420
rect 567896 52408 567902 52420
rect 579982 52408 579988 52420
rect 567896 52380 579988 52408
rect 567896 52368 567902 52380
rect 579982 52368 579988 52380
rect 580040 52368 580046 52420
rect 32490 52300 32496 52352
rect 32548 52340 32554 52352
rect 36722 52340 36728 52352
rect 32548 52312 36728 52340
rect 32548 52300 32554 52312
rect 36722 52300 36728 52312
rect 36780 52300 36786 52352
rect 29638 51620 29644 51672
rect 29696 51660 29702 51672
rect 34422 51660 34428 51672
rect 29696 51632 34428 51660
rect 29696 51620 29702 51632
rect 34422 51620 34428 51632
rect 34480 51620 34486 51672
rect 36814 51348 36820 51400
rect 36872 51388 36878 51400
rect 38102 51388 38108 51400
rect 36872 51360 38108 51388
rect 36872 51348 36878 51360
rect 38102 51348 38108 51360
rect 38160 51348 38166 51400
rect 41414 50844 41420 50856
rect 41375 50816 41420 50844
rect 41414 50804 41420 50816
rect 41472 50804 41478 50856
rect 40954 50668 40960 50720
rect 41012 50708 41018 50720
rect 41414 50708 41420 50720
rect 41012 50680 41420 50708
rect 41012 50668 41018 50680
rect 41414 50668 41420 50680
rect 41472 50668 41478 50720
rect 40310 50640 40316 50652
rect 40236 50612 40316 50640
rect 40236 50436 40264 50612
rect 40310 50600 40316 50612
rect 40368 50600 40374 50652
rect 40310 50464 40316 50516
rect 40368 50504 40374 50516
rect 40586 50504 40592 50516
rect 40368 50476 40592 50504
rect 40368 50464 40374 50476
rect 40586 50464 40592 50476
rect 40644 50464 40650 50516
rect 40236 50408 40540 50436
rect 40512 50312 40540 50408
rect 40494 50260 40500 50312
rect 40552 50260 40558 50312
rect 34514 49716 34520 49768
rect 34572 49756 34578 49768
rect 34572 49728 35894 49756
rect 34572 49716 34578 49728
rect 35866 49688 35894 49728
rect 38194 49688 38200 49700
rect 35866 49660 38200 49688
rect 38194 49648 38200 49660
rect 38252 49648 38258 49700
rect 2774 48288 2780 48340
rect 2832 48328 2838 48340
rect 4706 48328 4712 48340
rect 2832 48300 4712 48328
rect 2832 48288 2838 48300
rect 4706 48288 4712 48300
rect 4764 48288 4770 48340
rect 34514 47608 34520 47660
rect 34572 47648 34578 47660
rect 36262 47648 36268 47660
rect 34572 47620 36268 47648
rect 34572 47608 34578 47620
rect 36262 47608 36268 47620
rect 36320 47608 36326 47660
rect 559834 47472 559840 47524
rect 559892 47512 559898 47524
rect 564434 47512 564440 47524
rect 559892 47484 564440 47512
rect 559892 47472 559898 47484
rect 564434 47472 564440 47484
rect 564492 47472 564498 47524
rect 544654 46968 544660 46980
rect 544615 46940 544660 46968
rect 544654 46928 544660 46940
rect 544712 46928 544718 46980
rect 32398 46860 32404 46912
rect 32456 46900 32462 46912
rect 34514 46900 34520 46912
rect 32456 46872 34520 46900
rect 32456 46860 32462 46872
rect 34514 46860 34520 46872
rect 34572 46860 34578 46912
rect 36630 46860 36636 46912
rect 36688 46900 36694 46912
rect 37274 46900 37280 46912
rect 36688 46872 37280 46900
rect 36688 46860 36694 46872
rect 37274 46860 37280 46872
rect 37332 46860 37338 46912
rect 551554 46860 551560 46912
rect 551612 46900 551618 46912
rect 579982 46900 579988 46912
rect 551612 46872 579988 46900
rect 551612 46860 551618 46872
rect 579982 46860 579988 46872
rect 580040 46860 580046 46912
rect 544654 46792 544660 46844
rect 544712 46832 544718 46844
rect 563698 46832 563704 46844
rect 544712 46804 563704 46832
rect 544712 46792 544718 46804
rect 563698 46792 563704 46804
rect 563756 46792 563762 46844
rect 544654 46044 544660 46096
rect 544712 46084 544718 46096
rect 544838 46084 544844 46096
rect 544712 46056 544844 46084
rect 544712 46044 544718 46056
rect 544838 46044 544844 46056
rect 544896 46044 544902 46096
rect 544838 45908 544844 45960
rect 544896 45948 544902 45960
rect 545022 45948 545028 45960
rect 544896 45920 545028 45948
rect 544896 45908 544902 45920
rect 545022 45908 545028 45920
rect 545080 45908 545086 45960
rect 41782 45812 41788 45824
rect 41743 45784 41788 45812
rect 41782 45772 41788 45784
rect 41840 45772 41846 45824
rect 544657 45815 544715 45821
rect 544657 45781 544669 45815
rect 544703 45812 544715 45815
rect 545022 45812 545028 45824
rect 544703 45784 545028 45812
rect 544703 45781 544715 45784
rect 544657 45775 544715 45781
rect 545022 45772 545028 45784
rect 545080 45772 545086 45824
rect 41414 45704 41420 45756
rect 41472 45744 41478 45756
rect 41472 45716 41920 45744
rect 41472 45704 41478 45716
rect 40494 45568 40500 45620
rect 40552 45608 40558 45620
rect 40589 45611 40647 45617
rect 40589 45608 40601 45611
rect 40552 45580 40601 45608
rect 40552 45568 40558 45580
rect 40589 45577 40601 45580
rect 40635 45577 40647 45611
rect 41414 45608 41420 45620
rect 41375 45580 41420 45608
rect 40589 45571 40647 45577
rect 41414 45568 41420 45580
rect 41472 45568 41478 45620
rect 41892 45566 41920 45716
rect 559834 45608 559840 45620
rect 556172 45580 559840 45608
rect 41874 45514 41880 45566
rect 41932 45514 41938 45566
rect 552014 45500 552020 45552
rect 552072 45540 552078 45552
rect 556172 45540 556200 45580
rect 559834 45568 559840 45580
rect 559892 45568 559898 45620
rect 552072 45512 556200 45540
rect 552072 45500 552078 45512
rect 36262 44956 36268 45008
rect 36320 44996 36326 45008
rect 38838 44996 38844 45008
rect 36320 44968 38844 44996
rect 36320 44956 36326 44968
rect 38838 44956 38844 44968
rect 38896 44956 38902 45008
rect 3234 44752 3240 44804
rect 3292 44792 3298 44804
rect 3510 44792 3516 44804
rect 3292 44764 3516 44792
rect 3292 44752 3298 44764
rect 3510 44752 3516 44764
rect 3568 44752 3574 44804
rect 580534 44752 580540 44804
rect 580592 44792 580598 44804
rect 580718 44792 580724 44804
rect 580592 44764 580724 44792
rect 580592 44752 580598 44764
rect 580718 44752 580724 44764
rect 580776 44752 580782 44804
rect 37090 44616 37096 44668
rect 37148 44656 37154 44668
rect 41969 44659 42027 44665
rect 41969 44656 41981 44659
rect 37148 44628 41981 44656
rect 37148 44616 37154 44628
rect 41969 44625 41981 44628
rect 42015 44625 42027 44659
rect 542814 44656 542820 44668
rect 542775 44628 542820 44656
rect 41969 44619 42027 44625
rect 542814 44616 542820 44628
rect 542872 44616 542878 44668
rect 37550 44548 37556 44600
rect 37608 44588 37614 44600
rect 580902 44588 580908 44600
rect 37608 44560 580908 44588
rect 37608 44548 37614 44560
rect 580902 44548 580908 44560
rect 580960 44548 580966 44600
rect 3602 44480 3608 44532
rect 3660 44520 3666 44532
rect 3786 44520 3792 44532
rect 3660 44492 3792 44520
rect 3660 44480 3666 44492
rect 3786 44480 3792 44492
rect 3844 44480 3850 44532
rect 40586 44480 40592 44532
rect 40644 44520 40650 44532
rect 580074 44520 580080 44532
rect 40644 44492 580080 44520
rect 40644 44480 40650 44492
rect 580074 44480 580080 44492
rect 580132 44480 580138 44532
rect 38194 44412 38200 44464
rect 38252 44452 38258 44464
rect 38252 44424 40724 44452
rect 38252 44412 38258 44424
rect 40586 44384 40592 44396
rect 40547 44356 40592 44384
rect 40586 44344 40592 44356
rect 40644 44344 40650 44396
rect 40696 44384 40724 44424
rect 40954 44412 40960 44464
rect 41012 44452 41018 44464
rect 580442 44452 580448 44464
rect 41012 44424 580448 44452
rect 41012 44412 41018 44424
rect 580442 44412 580448 44424
rect 580500 44412 580506 44464
rect 41877 44387 41935 44393
rect 41877 44384 41889 44387
rect 40696 44356 41889 44384
rect 41877 44353 41889 44356
rect 41923 44353 41935 44387
rect 41877 44347 41935 44353
rect 41969 44387 42027 44393
rect 41969 44353 41981 44387
rect 42015 44384 42027 44387
rect 544930 44384 544936 44396
rect 42015 44356 544936 44384
rect 42015 44353 42027 44356
rect 41969 44347 42027 44353
rect 544930 44344 544936 44356
rect 544988 44344 544994 44396
rect 34422 44276 34428 44328
rect 34480 44316 34486 44328
rect 540977 44319 541035 44325
rect 540977 44316 540989 44319
rect 34480 44288 540989 44316
rect 34480 44276 34486 44288
rect 540977 44285 540989 44288
rect 541023 44285 541035 44319
rect 540977 44279 541035 44285
rect 541069 44319 541127 44325
rect 541069 44285 541081 44319
rect 541115 44316 541127 44319
rect 543642 44316 543648 44328
rect 541115 44288 543648 44316
rect 541115 44285 541127 44288
rect 541069 44279 541127 44285
rect 543642 44276 543648 44288
rect 543700 44276 543706 44328
rect 39206 44208 39212 44260
rect 39264 44248 39270 44260
rect 542170 44248 542176 44260
rect 39264 44220 542176 44248
rect 39264 44208 39270 44220
rect 542170 44208 542176 44220
rect 542228 44208 542234 44260
rect 542814 44208 542820 44260
rect 542872 44248 542878 44260
rect 544470 44248 544476 44260
rect 542872 44220 544476 44248
rect 542872 44208 542878 44220
rect 544470 44208 544476 44220
rect 544528 44208 544534 44260
rect 39022 44140 39028 44192
rect 39080 44180 39086 44192
rect 40954 44180 40960 44192
rect 39080 44152 40960 44180
rect 39080 44140 39086 44152
rect 40954 44140 40960 44152
rect 41012 44140 41018 44192
rect 41874 44180 41880 44192
rect 41835 44152 41880 44180
rect 41874 44140 41880 44152
rect 41932 44140 41938 44192
rect 542265 44183 542323 44189
rect 542265 44149 542277 44183
rect 542311 44180 542323 44183
rect 543366 44180 543372 44192
rect 542311 44152 543372 44180
rect 542311 44149 542323 44152
rect 542265 44143 542323 44149
rect 543366 44140 543372 44152
rect 543424 44140 543430 44192
rect 543550 44140 543556 44192
rect 543608 44180 543614 44192
rect 544746 44180 544752 44192
rect 543608 44152 544752 44180
rect 543608 44140 543614 44152
rect 544746 44140 544752 44152
rect 544804 44140 544810 44192
rect 34514 44072 34520 44124
rect 34572 44112 34578 44124
rect 544194 44112 544200 44124
rect 34572 44084 544200 44112
rect 34572 44072 34578 44084
rect 544194 44072 544200 44084
rect 544252 44072 544258 44124
rect 36538 44004 36544 44056
rect 36596 44044 36602 44056
rect 543918 44044 543924 44056
rect 36596 44016 543924 44044
rect 36596 44004 36602 44016
rect 543918 44004 543924 44016
rect 543976 44004 543982 44056
rect 39298 43936 39304 43988
rect 39356 43976 39362 43988
rect 39356 43948 542124 43976
rect 39356 43936 39362 43948
rect 39666 43868 39672 43920
rect 39724 43908 39730 43920
rect 542096 43908 542124 43948
rect 542170 43936 542176 43988
rect 542228 43976 542234 43988
rect 542265 43979 542323 43985
rect 542265 43976 542277 43979
rect 542228 43948 542277 43976
rect 542228 43936 542234 43948
rect 542265 43945 542277 43948
rect 542311 43945 542323 43979
rect 542265 43939 542323 43945
rect 546126 43908 546132 43920
rect 39724 43880 542032 43908
rect 542096 43880 546132 43908
rect 39724 43868 39730 43880
rect 38746 43800 38752 43852
rect 38804 43840 38810 43852
rect 541805 43843 541863 43849
rect 541805 43840 541817 43843
rect 38804 43812 541817 43840
rect 38804 43800 38810 43812
rect 541805 43809 541817 43812
rect 541851 43809 541863 43843
rect 542004 43840 542032 43880
rect 546126 43868 546132 43880
rect 546184 43868 546190 43920
rect 546402 43840 546408 43852
rect 542004 43812 546408 43840
rect 541805 43803 541863 43809
rect 546402 43800 546408 43812
rect 546460 43800 546466 43852
rect 39758 43732 39764 43784
rect 39816 43772 39822 43784
rect 546034 43772 546040 43784
rect 39816 43744 546040 43772
rect 39816 43732 39822 43744
rect 546034 43732 546040 43744
rect 546092 43732 546098 43784
rect 36722 43664 36728 43716
rect 36780 43704 36786 43716
rect 542722 43704 542728 43716
rect 36780 43676 542728 43704
rect 36780 43664 36786 43676
rect 542722 43664 542728 43676
rect 542780 43664 542786 43716
rect 41598 43596 41604 43648
rect 41656 43636 41662 43648
rect 541713 43639 541771 43645
rect 541713 43636 541725 43639
rect 41656 43608 541725 43636
rect 41656 43596 41662 43608
rect 541713 43605 541725 43608
rect 541759 43605 541771 43639
rect 541713 43599 541771 43605
rect 541805 43639 541863 43645
rect 541805 43605 541817 43639
rect 541851 43636 541863 43639
rect 546310 43636 546316 43648
rect 541851 43608 546316 43636
rect 541851 43605 541863 43608
rect 541805 43599 541863 43605
rect 546310 43596 546316 43608
rect 546368 43596 546374 43648
rect 37274 43528 37280 43580
rect 37332 43568 37338 43580
rect 541894 43568 541900 43580
rect 37332 43540 541900 43568
rect 37332 43528 37338 43540
rect 541894 43528 541900 43540
rect 541952 43528 541958 43580
rect 542722 43528 542728 43580
rect 542780 43568 542786 43580
rect 542817 43571 542875 43577
rect 542817 43568 542829 43571
rect 542780 43540 542829 43568
rect 542780 43528 542786 43540
rect 542817 43537 542829 43540
rect 542863 43537 542875 43571
rect 542817 43531 542875 43537
rect 20622 43460 20628 43512
rect 20680 43500 20686 43512
rect 544838 43500 544844 43512
rect 20680 43472 544844 43500
rect 20680 43460 20686 43472
rect 544838 43460 544844 43472
rect 544896 43460 544902 43512
rect 4798 43392 4804 43444
rect 4856 43432 4862 43444
rect 544286 43432 544292 43444
rect 4856 43404 544292 43432
rect 4856 43392 4862 43404
rect 544286 43392 544292 43404
rect 544344 43392 544350 43444
rect 41506 43324 41512 43376
rect 41564 43364 41570 43376
rect 544654 43364 544660 43376
rect 41564 43336 544660 43364
rect 41564 43324 41570 43336
rect 544654 43324 544660 43336
rect 544712 43324 544718 43376
rect 41874 43256 41880 43308
rect 41932 43296 41938 43308
rect 542814 43296 542820 43308
rect 41932 43268 542820 43296
rect 41932 43256 41938 43268
rect 542814 43256 542820 43268
rect 542872 43256 542878 43308
rect 41138 43188 41144 43240
rect 41196 43228 41202 43240
rect 542262 43228 542268 43240
rect 41196 43200 542268 43228
rect 41196 43188 41202 43200
rect 542262 43188 542268 43200
rect 542320 43188 542326 43240
rect 41322 43120 41328 43172
rect 41380 43160 41386 43172
rect 541069 43163 541127 43169
rect 541069 43160 541081 43163
rect 41380 43132 541081 43160
rect 41380 43120 41386 43132
rect 541069 43129 541081 43132
rect 541115 43129 541127 43163
rect 541069 43123 541127 43129
rect 541713 43163 541771 43169
rect 541713 43129 541725 43163
rect 541759 43160 541771 43163
rect 546218 43160 546224 43172
rect 541759 43132 546224 43160
rect 541759 43129 541771 43132
rect 541713 43123 541771 43129
rect 546218 43120 546224 43132
rect 546276 43120 546282 43172
rect 41414 43052 41420 43104
rect 41472 43092 41478 43104
rect 542170 43092 542176 43104
rect 41472 43064 542176 43092
rect 41472 43052 41478 43064
rect 542170 43052 542176 43064
rect 542228 43052 542234 43104
rect 41785 43027 41843 43033
rect 41785 42993 41797 43027
rect 41831 43024 41843 43027
rect 41874 43024 41880 43036
rect 41831 42996 41880 43024
rect 41831 42993 41843 42996
rect 41785 42987 41843 42993
rect 41874 42984 41880 42996
rect 41932 42984 41938 43036
rect 558178 42712 558184 42764
rect 558236 42752 558242 42764
rect 580166 42752 580172 42764
rect 558236 42724 580172 42752
rect 558236 42712 558242 42724
rect 580166 42712 580172 42724
rect 580224 42712 580230 42764
rect 536745 42619 536803 42625
rect 536745 42585 536757 42619
rect 536791 42616 536803 42619
rect 545298 42616 545304 42628
rect 536791 42588 545304 42616
rect 536791 42585 536803 42588
rect 536745 42579 536803 42585
rect 545298 42576 545304 42588
rect 545356 42576 545362 42628
rect 509145 42551 509203 42557
rect 509145 42517 509157 42551
rect 509191 42548 509203 42551
rect 543274 42548 543280 42560
rect 509191 42520 543280 42548
rect 509191 42517 509203 42520
rect 509145 42511 509203 42517
rect 543274 42508 543280 42520
rect 543332 42508 543338 42560
rect 40310 42440 40316 42492
rect 40368 42480 40374 42492
rect 191837 42483 191895 42489
rect 191837 42480 191849 42483
rect 40368 42452 191849 42480
rect 40368 42440 40374 42452
rect 191837 42449 191849 42452
rect 191883 42449 191895 42483
rect 191837 42443 191895 42449
rect 436005 42483 436063 42489
rect 436005 42449 436017 42483
rect 436051 42480 436063 42483
rect 543734 42480 543740 42492
rect 436051 42452 543740 42480
rect 436051 42449 436063 42452
rect 436005 42443 436063 42449
rect 543734 42440 543740 42452
rect 543792 42440 543798 42492
rect 40126 42372 40132 42424
rect 40184 42412 40190 42424
rect 196066 42412 196072 42424
rect 40184 42384 196072 42412
rect 40184 42372 40190 42384
rect 196066 42372 196072 42384
rect 196124 42372 196130 42424
rect 379422 42372 379428 42424
rect 379480 42412 379486 42424
rect 542446 42412 542452 42424
rect 379480 42384 542452 42412
rect 379480 42372 379486 42384
rect 542446 42372 542452 42384
rect 542504 42372 542510 42424
rect 38930 42304 38936 42356
rect 38988 42344 38994 42356
rect 231854 42344 231860 42356
rect 38988 42316 231860 42344
rect 38988 42304 38994 42316
rect 231854 42304 231860 42316
rect 231912 42304 231918 42356
rect 277302 42304 277308 42356
rect 277360 42344 277366 42356
rect 545022 42344 545028 42356
rect 277360 42316 545028 42344
rect 277360 42304 277366 42316
rect 545022 42304 545028 42316
rect 545080 42304 545086 42356
rect 4154 42236 4160 42288
rect 4212 42276 4218 42288
rect 320174 42276 320180 42288
rect 4212 42248 320180 42276
rect 4212 42236 4218 42248
rect 320174 42236 320180 42248
rect 320232 42236 320238 42288
rect 333882 42236 333888 42288
rect 333940 42276 333946 42288
rect 543826 42276 543832 42288
rect 333940 42248 543832 42276
rect 333940 42236 333946 42248
rect 543826 42236 543832 42248
rect 543884 42236 543890 42288
rect 40586 42168 40592 42220
rect 40644 42208 40650 42220
rect 382274 42208 382280 42220
rect 40644 42180 382280 42208
rect 40644 42168 40650 42180
rect 382274 42168 382280 42180
rect 382332 42168 382338 42220
rect 395982 42168 395988 42220
rect 396040 42208 396046 42220
rect 543458 42208 543464 42220
rect 396040 42180 543464 42208
rect 396040 42168 396046 42180
rect 543458 42168 543464 42180
rect 543516 42168 543522 42220
rect 169662 42100 169668 42152
rect 169720 42140 169726 42152
rect 544378 42140 544384 42152
rect 169720 42112 544384 42140
rect 169720 42100 169726 42112
rect 544378 42100 544384 42112
rect 544436 42100 544442 42152
rect 39942 42032 39948 42084
rect 40000 42072 40006 42084
rect 580442 42072 580448 42084
rect 40000 42044 580448 42072
rect 40000 42032 40006 42044
rect 580442 42032 580448 42044
rect 580500 42032 580506 42084
rect 191834 42004 191840 42016
rect 191795 41976 191840 42004
rect 191834 41964 191840 41976
rect 191892 41964 191898 42016
rect 436002 42004 436008 42016
rect 435963 41976 436008 42004
rect 436002 41964 436008 41976
rect 436060 41964 436066 42016
rect 509142 42004 509148 42016
rect 509103 41976 509148 42004
rect 509142 41964 509148 41976
rect 509200 41964 509206 42016
rect 536742 42004 536748 42016
rect 536703 41976 536748 42004
rect 536742 41964 536748 41976
rect 536800 41964 536806 42016
rect 538306 41420 538312 41472
rect 538364 41460 538370 41472
rect 542354 41460 542360 41472
rect 538364 41432 542360 41460
rect 538364 41420 538370 41432
rect 542354 41420 542360 41432
rect 542412 41420 542418 41472
rect 3326 41352 3332 41404
rect 3384 41392 3390 41404
rect 65978 41392 65984 41404
rect 3384 41364 65984 41392
rect 3384 41352 3390 41364
rect 65978 41352 65984 41364
rect 66036 41352 66042 41404
rect 157426 41352 157432 41404
rect 157484 41392 157490 41404
rect 162854 41392 162860 41404
rect 157484 41364 162860 41392
rect 157484 41352 157490 41364
rect 162854 41352 162860 41364
rect 162912 41352 162918 41404
rect 384666 41352 384672 41404
rect 384724 41392 384730 41404
rect 547690 41392 547696 41404
rect 384724 41364 547696 41392
rect 384724 41352 384730 41364
rect 547690 41352 547696 41364
rect 547748 41352 547754 41404
rect 7834 41284 7840 41336
rect 7892 41324 7898 41336
rect 71774 41324 71780 41336
rect 7892 41296 71780 41324
rect 7892 41284 7898 41296
rect 71774 41284 71780 41296
rect 71832 41284 71838 41336
rect 305914 41284 305920 41336
rect 305972 41324 305978 41336
rect 547782 41324 547788 41336
rect 305972 41296 547788 41324
rect 305972 41284 305978 41296
rect 547782 41284 547788 41296
rect 547840 41284 547846 41336
rect 7558 41216 7564 41268
rect 7616 41256 7622 41268
rect 156598 41256 156604 41268
rect 7616 41228 156604 41256
rect 7616 41216 7622 41228
rect 156598 41216 156604 41228
rect 156656 41216 156662 41268
rect 275554 41216 275560 41268
rect 275612 41256 275618 41268
rect 547230 41256 547236 41268
rect 275612 41228 547236 41256
rect 275612 41216 275618 41228
rect 547230 41216 547236 41228
rect 547288 41216 547294 41268
rect 33042 41148 33048 41200
rect 33100 41188 33106 41200
rect 329190 41188 329196 41200
rect 33100 41160 329196 41188
rect 33100 41148 33106 41160
rect 329190 41148 329196 41160
rect 329248 41148 329254 41200
rect 366450 41148 366456 41200
rect 366508 41188 366514 41200
rect 552750 41188 552756 41200
rect 366508 41160 552756 41188
rect 366508 41148 366514 41160
rect 552750 41148 552756 41160
rect 552808 41148 552814 41200
rect 9122 41080 9128 41132
rect 9180 41120 9186 41132
rect 168742 41120 168748 41132
rect 9180 41092 168748 41120
rect 9180 41080 9186 41092
rect 168742 41080 168748 41092
rect 168800 41080 168806 41132
rect 245194 41080 245200 41132
rect 245252 41120 245258 41132
rect 548518 41120 548524 41132
rect 245252 41092 548524 41120
rect 245252 41080 245258 41092
rect 548518 41080 548524 41092
rect 548576 41080 548582 41132
rect 5258 41012 5264 41064
rect 5316 41052 5322 41064
rect 226334 41052 226340 41064
rect 5316 41024 226340 41052
rect 5316 41012 5322 41024
rect 226334 41012 226340 41024
rect 226392 41012 226398 41064
rect 269482 41012 269488 41064
rect 269540 41052 269546 41064
rect 580350 41052 580356 41064
rect 269540 41024 580356 41052
rect 269540 41012 269546 41024
rect 580350 41012 580356 41024
rect 580408 41012 580414 41064
rect 4890 40944 4896 40996
rect 4948 40984 4954 40996
rect 232774 40984 232780 40996
rect 4948 40956 232780 40984
rect 4948 40944 4954 40956
rect 232774 40944 232780 40956
rect 232832 40944 232838 40996
rect 238754 40944 238760 40996
rect 238812 40984 238818 40996
rect 571334 40984 571340 40996
rect 238812 40956 571340 40984
rect 238812 40944 238818 40956
rect 571334 40944 571340 40956
rect 571392 40944 571398 40996
rect 7742 40876 7748 40928
rect 7800 40916 7806 40928
rect 347774 40916 347780 40928
rect 7800 40888 347780 40916
rect 7800 40876 7806 40888
rect 347774 40876 347780 40888
rect 347832 40876 347838 40928
rect 350994 40876 351000 40928
rect 351052 40916 351058 40928
rect 548978 40916 548984 40928
rect 351052 40888 548984 40916
rect 351052 40876 351058 40888
rect 548978 40876 548984 40888
rect 549036 40876 549042 40928
rect 6546 40808 6552 40860
rect 6604 40848 6610 40860
rect 408310 40848 408316 40860
rect 6604 40820 408316 40848
rect 6604 40808 6610 40820
rect 408310 40808 408316 40820
rect 408368 40808 408374 40860
rect 3418 40740 3424 40792
rect 3476 40780 3482 40792
rect 411438 40780 411444 40792
rect 3476 40752 411444 40780
rect 3476 40740 3482 40752
rect 411438 40740 411444 40752
rect 411496 40740 411502 40792
rect 5350 40672 5356 40724
rect 5408 40712 5414 40724
rect 420454 40712 420460 40724
rect 5408 40684 420460 40712
rect 5408 40672 5414 40684
rect 420454 40672 420460 40684
rect 420512 40672 420518 40724
rect 513282 40672 513288 40724
rect 513340 40712 513346 40724
rect 542722 40712 542728 40724
rect 513340 40684 542728 40712
rect 513340 40672 513346 40684
rect 542722 40672 542728 40684
rect 542780 40672 542786 40724
rect 4706 40604 4712 40656
rect 4764 40644 4770 40656
rect 69198 40644 69204 40656
rect 4764 40616 69204 40644
rect 4764 40604 4770 40616
rect 69198 40604 69204 40616
rect 69256 40604 69262 40656
rect 150986 40604 150992 40656
rect 151044 40644 151050 40656
rect 580810 40644 580816 40656
rect 151044 40616 580816 40644
rect 151044 40604 151050 40616
rect 580810 40604 580816 40616
rect 580868 40604 580874 40656
rect 9030 40536 9036 40588
rect 9088 40576 9094 40588
rect 441614 40576 441620 40588
rect 9088 40548 441620 40576
rect 9088 40536 9094 40548
rect 441614 40536 441620 40548
rect 441672 40536 441678 40588
rect 493226 40536 493232 40588
rect 493284 40576 493290 40588
rect 545850 40576 545856 40588
rect 493284 40548 545856 40576
rect 493284 40536 493290 40548
rect 545850 40536 545856 40548
rect 545908 40536 545914 40588
rect 68002 40468 68008 40520
rect 68060 40508 68066 40520
rect 135806 40508 135812 40520
rect 68060 40480 135812 40508
rect 68060 40468 68066 40480
rect 135806 40468 135812 40480
rect 135864 40468 135870 40520
rect 138842 40468 138848 40520
rect 138900 40508 138906 40520
rect 580626 40508 580632 40520
rect 138900 40480 580632 40508
rect 138900 40468 138906 40480
rect 580626 40468 580632 40480
rect 580684 40468 580690 40520
rect 7926 40400 7932 40452
rect 7984 40440 7990 40452
rect 96430 40440 96436 40452
rect 7984 40412 96436 40440
rect 7984 40400 7990 40412
rect 96430 40400 96436 40412
rect 96488 40400 96494 40452
rect 102594 40400 102600 40452
rect 102652 40440 102658 40452
rect 547506 40440 547512 40452
rect 102652 40412 547512 40440
rect 102652 40400 102658 40412
rect 547506 40400 547512 40412
rect 547564 40400 547570 40452
rect 3970 40332 3976 40384
rect 4028 40372 4034 40384
rect 465902 40372 465908 40384
rect 4028 40344 465908 40372
rect 4028 40332 4034 40344
rect 465902 40332 465908 40344
rect 465960 40332 465966 40384
rect 469122 40332 469128 40384
rect 469180 40372 469186 40384
rect 580074 40372 580080 40384
rect 469180 40344 580080 40372
rect 469180 40332 469186 40344
rect 580074 40332 580080 40344
rect 580132 40332 580138 40384
rect 5074 40264 5080 40316
rect 5132 40304 5138 40316
rect 474918 40304 474924 40316
rect 5132 40276 474924 40304
rect 5132 40264 5138 40276
rect 474918 40264 474924 40276
rect 474976 40264 474982 40316
rect 496354 40264 496360 40316
rect 496412 40304 496418 40316
rect 580534 40304 580540 40316
rect 496412 40276 580540 40304
rect 496412 40264 496418 40276
rect 580534 40264 580540 40276
rect 580592 40264 580598 40316
rect 5442 40196 5448 40248
rect 5500 40236 5506 40248
rect 499206 40236 499212 40248
rect 5500 40208 499212 40236
rect 5500 40196 5506 40208
rect 499206 40196 499212 40208
rect 499264 40196 499270 40248
rect 3786 40128 3792 40180
rect 3844 40168 3850 40180
rect 508406 40168 508412 40180
rect 3844 40140 508412 40168
rect 3844 40128 3850 40140
rect 508406 40128 508412 40140
rect 508464 40128 508470 40180
rect 6730 40060 6736 40112
rect 6788 40100 6794 40112
rect 520366 40100 520372 40112
rect 6788 40072 520372 40100
rect 6788 40060 6794 40072
rect 520366 40060 520372 40072
rect 520424 40060 520430 40112
rect 37182 39992 37188 40044
rect 37240 40032 37246 40044
rect 51074 40032 51080 40044
rect 37240 40004 51080 40032
rect 37240 39992 37246 40004
rect 51074 39992 51080 40004
rect 51132 39992 51138 40044
rect 123754 39992 123760 40044
rect 123812 40032 123818 40044
rect 131117 40035 131175 40041
rect 131117 40032 131129 40035
rect 123812 40004 131129 40032
rect 123812 39992 123818 40004
rect 131117 40001 131129 40004
rect 131163 40001 131175 40035
rect 131117 39995 131175 40001
rect 345658 39992 345664 40044
rect 345716 40032 345722 40044
rect 348234 40032 348240 40044
rect 345716 40004 348240 40032
rect 345716 39992 345722 40004
rect 348234 39992 348240 40004
rect 348292 39992 348298 40044
rect 352374 39992 352380 40044
rect 352432 40032 352438 40044
rect 354950 40032 354956 40044
rect 352432 40004 354956 40032
rect 352432 39992 352438 40004
rect 354950 39992 354956 40004
rect 355008 39992 355014 40044
rect 511442 39992 511448 40044
rect 511500 40032 511506 40044
rect 548886 40032 548892 40044
rect 511500 40004 548892 40032
rect 511500 39992 511506 40004
rect 548886 39992 548892 40004
rect 548944 39992 548950 40044
rect 41782 39924 41788 39976
rect 41840 39964 41846 39976
rect 159910 39964 159916 39976
rect 41840 39936 159916 39964
rect 41840 39924 41846 39936
rect 159910 39924 159916 39936
rect 159968 39924 159974 39976
rect 314562 39924 314568 39976
rect 314620 39964 314626 39976
rect 316034 39964 316040 39976
rect 314620 39936 316040 39964
rect 314620 39924 314626 39936
rect 316034 39924 316040 39936
rect 316092 39924 316098 39976
rect 529658 39924 529664 39976
rect 529716 39964 529722 39976
rect 552934 39964 552940 39976
rect 529716 39936 552940 39964
rect 529716 39924 529722 39936
rect 552934 39924 552940 39936
rect 552992 39924 552998 39976
rect 5166 39856 5172 39908
rect 5224 39896 5230 39908
rect 429654 39896 429660 39908
rect 5224 39868 429660 39896
rect 5224 39856 5230 39868
rect 429654 39856 429660 39868
rect 429712 39856 429718 39908
rect 535730 39856 535736 39908
rect 535788 39896 535794 39908
rect 551462 39896 551468 39908
rect 535788 39868 551468 39896
rect 535788 39856 535794 39868
rect 551462 39856 551468 39868
rect 551520 39856 551526 39908
rect 3602 39788 3608 39840
rect 3660 39828 3666 39840
rect 417510 39828 417516 39840
rect 3660 39800 417516 39828
rect 3660 39788 3666 39800
rect 417510 39788 417516 39800
rect 417568 39788 417574 39840
rect 426618 39788 426624 39840
rect 426676 39828 426682 39840
rect 439498 39828 439504 39840
rect 426676 39800 439504 39828
rect 426676 39788 426682 39800
rect 439498 39788 439504 39800
rect 439556 39788 439562 39840
rect 450906 39788 450912 39840
rect 450964 39828 450970 39840
rect 548794 39828 548800 39840
rect 450964 39800 548800 39828
rect 450964 39788 450970 39800
rect 548794 39788 548800 39800
rect 548852 39788 548858 39840
rect 1302 39720 1308 39772
rect 1360 39760 1366 39772
rect 41966 39760 41972 39772
rect 1360 39732 41972 39760
rect 1360 39720 1366 39732
rect 41966 39720 41972 39732
rect 42024 39720 42030 39772
rect 65978 39720 65984 39772
rect 66036 39760 66042 39772
rect 453758 39760 453764 39772
rect 66036 39732 453764 39760
rect 66036 39720 66042 39732
rect 453758 39720 453764 39732
rect 453816 39720 453822 39772
rect 459922 39720 459928 39772
rect 459980 39760 459986 39772
rect 547598 39760 547604 39772
rect 459980 39732 547604 39760
rect 459980 39720 459986 39732
rect 547598 39720 547604 39732
rect 547656 39720 547662 39772
rect 2774 39652 2780 39704
rect 2832 39692 2838 39704
rect 4982 39692 4988 39704
rect 2832 39664 4988 39692
rect 2832 39652 2838 39664
rect 4982 39652 4988 39664
rect 5040 39652 5046 39704
rect 9490 39652 9496 39704
rect 9548 39692 9554 39704
rect 196342 39692 196348 39704
rect 9548 39664 196348 39692
rect 9548 39652 9554 39664
rect 196342 39652 196348 39664
rect 196400 39652 196406 39704
rect 208578 39652 208584 39704
rect 208636 39692 208642 39704
rect 551922 39692 551928 39704
rect 208636 39664 551928 39692
rect 208636 39652 208642 39664
rect 551922 39652 551928 39664
rect 551980 39652 551986 39704
rect 9214 39584 9220 39636
rect 9272 39624 9278 39636
rect 190270 39624 190276 39636
rect 9272 39596 190276 39624
rect 9272 39584 9278 39596
rect 190270 39584 190276 39596
rect 190328 39584 190334 39636
rect 211522 39584 211528 39636
rect 211580 39624 211586 39636
rect 549070 39624 549076 39636
rect 211580 39596 549076 39624
rect 211580 39584 211586 39596
rect 549070 39584 549076 39596
rect 549128 39584 549134 39636
rect 8202 39516 8208 39568
rect 8260 39556 8266 39568
rect 214558 39556 214564 39568
rect 8260 39528 214564 39556
rect 8260 39516 8266 39528
rect 214558 39516 214564 39528
rect 214616 39516 214622 39568
rect 217594 39516 217600 39568
rect 217652 39556 217658 39568
rect 550358 39556 550364 39568
rect 217652 39528 550364 39556
rect 217652 39516 217658 39528
rect 550358 39516 550364 39528
rect 550416 39516 550422 39568
rect 9306 39448 9312 39500
rect 9364 39488 9370 39500
rect 338758 39488 338764 39500
rect 9364 39460 338764 39488
rect 9364 39448 9370 39460
rect 338758 39448 338764 39460
rect 338816 39448 338822 39500
rect 344922 39448 344928 39500
rect 344980 39488 344986 39500
rect 542909 39491 542967 39497
rect 542909 39488 542921 39491
rect 344980 39460 542921 39488
rect 344980 39448 344986 39460
rect 542909 39457 542921 39460
rect 542955 39457 542967 39491
rect 542909 39451 542967 39457
rect 543001 39491 543059 39497
rect 543001 39457 543013 39491
rect 543047 39488 543059 39491
rect 550082 39488 550088 39500
rect 543047 39460 550088 39488
rect 543047 39457 543059 39460
rect 543001 39451 543059 39457
rect 550082 39448 550088 39460
rect 550140 39448 550146 39500
rect 8110 39380 8116 39432
rect 8168 39420 8174 39432
rect 335630 39420 335636 39432
rect 8168 39392 335636 39420
rect 8168 39380 8174 39392
rect 335630 39380 335636 39392
rect 335688 39380 335694 39432
rect 369026 39380 369032 39432
rect 369084 39420 369090 39432
rect 551738 39420 551744 39432
rect 369084 39392 551744 39420
rect 369084 39380 369090 39392
rect 551738 39380 551744 39392
rect 551796 39380 551802 39432
rect 13722 39312 13728 39364
rect 13780 39352 13786 39364
rect 53926 39352 53932 39364
rect 13780 39324 53932 39352
rect 13780 39312 13786 39324
rect 53926 39312 53932 39324
rect 53984 39312 53990 39364
rect 59354 39312 59360 39364
rect 59412 39352 59418 39364
rect 61378 39352 61384 39364
rect 59412 39324 61384 39352
rect 59412 39312 59418 39324
rect 61378 39312 61384 39324
rect 61436 39312 61442 39364
rect 86862 39312 86868 39364
rect 86920 39352 86926 39364
rect 117590 39352 117596 39364
rect 86920 39324 117596 39352
rect 86920 39312 86926 39324
rect 117590 39312 117596 39324
rect 117648 39312 117654 39364
rect 126698 39312 126704 39364
rect 126756 39352 126762 39364
rect 443638 39352 443644 39364
rect 126756 39324 443644 39352
rect 126756 39312 126762 39324
rect 443638 39312 443644 39324
rect 443696 39312 443702 39364
rect 514386 39312 514392 39364
rect 514444 39352 514450 39364
rect 580258 39352 580264 39364
rect 514444 39324 580264 39352
rect 514444 39312 514450 39324
rect 580258 39312 580264 39324
rect 580316 39312 580322 39364
rect 6086 39244 6092 39296
rect 6144 39284 6150 39296
rect 302326 39284 302332 39296
rect 6144 39256 302332 39284
rect 6144 39244 6150 39256
rect 302326 39244 302332 39256
rect 302384 39244 302390 39296
rect 332778 39244 332784 39296
rect 332836 39284 332842 39296
rect 367738 39284 367744 39296
rect 332836 39256 367744 39284
rect 332836 39244 332842 39256
rect 367738 39244 367744 39256
rect 367796 39244 367802 39296
rect 375098 39244 375104 39296
rect 375156 39284 375162 39296
rect 385034 39284 385040 39296
rect 375156 39256 385040 39284
rect 375156 39244 375162 39256
rect 385034 39244 385040 39256
rect 385092 39244 385098 39296
rect 387242 39244 387248 39296
rect 387300 39284 387306 39296
rect 549898 39284 549904 39296
rect 387300 39256 549904 39284
rect 387300 39244 387306 39256
rect 549898 39244 549904 39256
rect 549956 39244 549962 39296
rect 9398 39176 9404 39228
rect 9456 39216 9462 39228
rect 250806 39216 250812 39228
rect 9456 39188 250812 39216
rect 9456 39176 9462 39188
rect 250806 39176 250812 39188
rect 250864 39176 250870 39228
rect 260098 39176 260104 39228
rect 260156 39216 260162 39228
rect 543001 39219 543059 39225
rect 543001 39216 543013 39219
rect 260156 39188 543013 39216
rect 260156 39176 260162 39188
rect 543001 39185 543013 39188
rect 543047 39185 543059 39219
rect 543001 39179 543059 39185
rect 10870 39108 10876 39160
rect 10928 39148 10934 39160
rect 241790 39148 241796 39160
rect 10928 39120 241796 39148
rect 10928 39108 10934 39120
rect 241790 39108 241796 39120
rect 241848 39108 241854 39160
rect 247954 39108 247960 39160
rect 248012 39148 248018 39160
rect 259454 39148 259460 39160
rect 248012 39120 259460 39148
rect 248012 39108 248018 39120
rect 259454 39108 259460 39120
rect 259512 39108 259518 39160
rect 281258 39108 281264 39160
rect 281316 39148 281322 39160
rect 551830 39148 551836 39160
rect 281316 39120 551836 39148
rect 281316 39108 281322 39120
rect 551830 39108 551836 39120
rect 551888 39108 551894 39160
rect 3510 39040 3516 39092
rect 3568 39080 3574 39092
rect 178126 39080 178132 39092
rect 3568 39052 178132 39080
rect 3568 39040 3574 39052
rect 178126 39040 178132 39052
rect 178184 39040 178190 39092
rect 205450 39040 205456 39092
rect 205508 39080 205514 39092
rect 285674 39080 285680 39092
rect 205508 39052 285680 39080
rect 205508 39040 205514 39052
rect 285674 39040 285680 39052
rect 285732 39040 285738 39092
rect 290274 39040 290280 39092
rect 290332 39080 290338 39092
rect 548610 39080 548616 39092
rect 290332 39052 548616 39080
rect 290332 39040 290338 39052
rect 548610 39040 548616 39052
rect 548668 39040 548674 39092
rect 38378 38972 38384 39024
rect 38436 39012 38442 39024
rect 181254 39012 181260 39024
rect 38436 38984 181260 39012
rect 38436 38972 38442 38984
rect 181254 38972 181260 38984
rect 181312 38972 181318 39024
rect 272242 38972 272248 39024
rect 272300 39012 272306 39024
rect 301498 39012 301504 39024
rect 272300 38984 301504 39012
rect 272300 38972 272306 38984
rect 301498 38972 301504 38984
rect 301556 38972 301562 39024
rect 362954 38972 362960 39024
rect 363012 39012 363018 39024
rect 372614 39012 372620 39024
rect 363012 38984 372620 39012
rect 363012 38972 363018 38984
rect 372614 38972 372620 38984
rect 372672 38972 372678 39024
rect 435634 38972 435640 39024
rect 435692 39012 435698 39024
rect 451918 39012 451924 39024
rect 435692 38984 451924 39012
rect 435692 38972 435698 38984
rect 451918 38972 451924 38984
rect 451976 38972 451982 39024
rect 490282 38972 490288 39024
rect 490340 39012 490346 39024
rect 548702 39012 548708 39024
rect 490340 38984 548708 39012
rect 490340 38972 490346 38984
rect 548702 38972 548708 38984
rect 548760 38972 548766 39024
rect 44082 38904 44088 38956
rect 44140 38944 44146 38956
rect 81158 38944 81164 38956
rect 44140 38916 81164 38944
rect 44140 38904 44146 38916
rect 81158 38904 81164 38916
rect 81216 38904 81222 38956
rect 105538 38904 105544 38956
rect 105596 38944 105602 38956
rect 159358 38944 159364 38956
rect 105596 38916 159364 38944
rect 105596 38904 105602 38916
rect 159358 38904 159364 38916
rect 159416 38904 159422 38956
rect 266262 38904 266268 38956
rect 266320 38944 266326 38956
rect 293310 38944 293316 38956
rect 266320 38916 293316 38944
rect 266320 38904 266326 38916
rect 293310 38904 293316 38916
rect 293368 38904 293374 38956
rect 502426 38904 502432 38956
rect 502484 38944 502490 38956
rect 547874 38944 547880 38956
rect 502484 38916 547880 38944
rect 502484 38904 502490 38916
rect 547874 38904 547880 38916
rect 547932 38904 547938 38956
rect 38286 38836 38292 38888
rect 38344 38876 38350 38888
rect 47854 38876 47860 38888
rect 38344 38848 47860 38876
rect 38344 38836 38350 38848
rect 47854 38836 47860 38848
rect 47912 38836 47918 38888
rect 90450 38836 90456 38888
rect 90508 38876 90514 38888
rect 131758 38876 131764 38888
rect 90508 38848 131764 38876
rect 90508 38836 90514 38848
rect 131758 38836 131764 38848
rect 131816 38836 131822 38888
rect 131850 38836 131856 38888
rect 131908 38876 131914 38888
rect 172054 38876 172060 38888
rect 131908 38848 172060 38876
rect 131908 38836 131914 38848
rect 172054 38836 172060 38848
rect 172112 38836 172118 38888
rect 444834 38836 444840 38888
rect 444892 38876 444898 38888
rect 444892 38848 541756 38876
rect 444892 38836 444898 38848
rect 6454 38768 6460 38820
rect 6512 38808 6518 38820
rect 114646 38808 114652 38820
rect 6512 38780 114652 38808
rect 6512 38768 6518 38780
rect 114646 38768 114652 38780
rect 114704 38768 114710 38820
rect 119982 38768 119988 38820
rect 120040 38808 120046 38820
rect 144914 38808 144920 38820
rect 120040 38780 144920 38808
rect 120040 38768 120046 38780
rect 144914 38768 144920 38780
rect 144972 38768 144978 38820
rect 154114 38768 154120 38820
rect 154172 38808 154178 38820
rect 182818 38808 182824 38820
rect 154172 38780 182824 38808
rect 154172 38768 154178 38780
rect 182818 38768 182824 38780
rect 182876 38768 182882 38820
rect 254026 38768 254032 38820
rect 254084 38808 254090 38820
rect 255222 38808 255228 38820
rect 254084 38780 255228 38808
rect 254084 38768 254090 38780
rect 255222 38768 255228 38780
rect 255280 38768 255286 38820
rect 414474 38768 414480 38820
rect 414532 38808 414538 38820
rect 415302 38808 415308 38820
rect 414532 38780 415308 38808
rect 414532 38768 414538 38780
rect 415302 38768 415308 38780
rect 415360 38768 415366 38820
rect 482922 38768 482928 38820
rect 482980 38808 482986 38820
rect 484118 38808 484124 38820
rect 482980 38780 484124 38808
rect 482980 38768 482986 38780
rect 484118 38768 484124 38780
rect 484176 38768 484182 38820
rect 538674 38768 538680 38820
rect 538732 38808 538738 38820
rect 539502 38808 539508 38820
rect 538732 38780 539508 38808
rect 538732 38768 538738 38780
rect 539502 38768 539508 38780
rect 539560 38768 539566 38820
rect 541728 38808 541756 38848
rect 541802 38836 541808 38888
rect 541860 38876 541866 38888
rect 542262 38876 542268 38888
rect 541860 38848 542268 38876
rect 541860 38836 541866 38848
rect 542262 38836 542268 38848
rect 542320 38836 542326 38888
rect 542909 38879 542967 38885
rect 542909 38845 542921 38879
rect 542955 38876 542967 38879
rect 550542 38876 550548 38888
rect 542955 38848 550548 38876
rect 542955 38845 542967 38848
rect 542909 38839 542967 38845
rect 550542 38836 550548 38848
rect 550600 38836 550606 38888
rect 550174 38808 550180 38820
rect 541728 38780 550180 38808
rect 550174 38768 550180 38780
rect 550232 38768 550238 38820
rect 41874 38700 41880 38752
rect 41932 38740 41938 38752
rect 75270 38740 75276 38752
rect 41932 38712 75276 38740
rect 41932 38700 41938 38712
rect 75270 38700 75276 38712
rect 75328 38700 75334 38752
rect 129826 38700 129832 38752
rect 129884 38740 129890 38752
rect 131022 38740 131028 38752
rect 129884 38712 131028 38740
rect 129884 38700 129890 38712
rect 131022 38700 131028 38712
rect 131080 38700 131086 38752
rect 131117 38743 131175 38749
rect 131117 38709 131129 38743
rect 131163 38740 131175 38743
rect 550266 38740 550272 38752
rect 131163 38712 550272 38740
rect 131163 38709 131175 38712
rect 131117 38703 131175 38709
rect 550266 38700 550272 38712
rect 550324 38700 550330 38752
rect 7650 38632 7656 38684
rect 7708 38672 7714 38684
rect 44910 38672 44916 38684
rect 7708 38644 44916 38672
rect 7708 38632 7714 38644
rect 44910 38632 44916 38644
rect 44968 38632 44974 38684
rect 108666 38632 108672 38684
rect 108724 38672 108730 38684
rect 552842 38672 552848 38684
rect 108724 38644 552848 38672
rect 108724 38632 108730 38644
rect 552842 38632 552848 38644
rect 552900 38632 552906 38684
rect 346302 38292 346308 38344
rect 346360 38332 346366 38344
rect 350534 38332 350540 38344
rect 346360 38304 350540 38332
rect 346360 38292 346366 38304
rect 350534 38292 350540 38304
rect 350592 38292 350598 38344
rect 349982 37884 349988 37936
rect 350040 37924 350046 37936
rect 352374 37924 352380 37936
rect 350040 37896 352380 37924
rect 350040 37884 350046 37896
rect 352374 37884 352380 37896
rect 352432 37884 352438 37936
rect 449802 37884 449808 37936
rect 449860 37924 449866 37936
rect 544562 37924 544568 37936
rect 449860 37896 544568 37924
rect 449860 37884 449866 37896
rect 544562 37884 544568 37896
rect 544620 37884 544626 37936
rect 547138 37204 547144 37256
rect 547196 37244 547202 37256
rect 580166 37244 580172 37256
rect 547196 37216 580172 37244
rect 547196 37204 547202 37216
rect 580166 37204 580172 37216
rect 580224 37204 580230 37256
rect 39482 36524 39488 36576
rect 39540 36564 39546 36576
rect 368474 36564 368480 36576
rect 39540 36536 368480 36564
rect 39540 36524 39546 36536
rect 368474 36524 368480 36536
rect 368532 36524 368538 36576
rect 343542 35912 343548 35964
rect 343600 35952 343606 35964
rect 346302 35952 346308 35964
rect 343600 35924 346308 35952
rect 343600 35912 343606 35924
rect 346302 35912 346308 35924
rect 346360 35912 346366 35964
rect 343634 35232 343640 35284
rect 343692 35272 343698 35284
rect 349982 35272 349988 35284
rect 343692 35244 349988 35272
rect 343692 35232 343698 35244
rect 349982 35232 349988 35244
rect 350040 35232 350046 35284
rect 40034 35164 40040 35216
rect 40092 35204 40098 35216
rect 349154 35204 349160 35216
rect 40092 35176 349160 35204
rect 40092 35164 40098 35176
rect 349154 35164 349160 35176
rect 349212 35164 349218 35216
rect 345658 34524 345664 34536
rect 344986 34496 345664 34524
rect 340506 34416 340512 34468
rect 340564 34456 340570 34468
rect 344986 34456 345014 34496
rect 345658 34484 345664 34496
rect 345716 34484 345722 34536
rect 340564 34428 345014 34456
rect 340564 34416 340570 34428
rect 3418 34348 3424 34400
rect 3476 34388 3482 34400
rect 8938 34388 8944 34400
rect 3476 34360 8944 34388
rect 3476 34348 3482 34360
rect 8938 34348 8944 34360
rect 8996 34348 9002 34400
rect 341518 33124 341524 33176
rect 341576 33164 341582 33176
rect 343542 33164 343548 33176
rect 341576 33136 343548 33164
rect 341576 33124 341582 33136
rect 343542 33124 343548 33136
rect 343600 33124 343606 33176
rect 438762 33056 438768 33108
rect 438820 33096 438826 33108
rect 580074 33096 580080 33108
rect 438820 33068 580080 33096
rect 438820 33056 438826 33068
rect 580074 33056 580080 33068
rect 580132 33056 580138 33108
rect 340506 31804 340512 31816
rect 338132 31776 340512 31804
rect 335998 31696 336004 31748
rect 336056 31736 336062 31748
rect 338132 31736 338160 31776
rect 340506 31764 340512 31776
rect 340564 31764 340570 31816
rect 343634 31804 343640 31816
rect 340892 31776 343640 31804
rect 336056 31708 338160 31736
rect 336056 31696 336062 31708
rect 339678 31696 339684 31748
rect 339736 31736 339742 31748
rect 340892 31736 340920 31776
rect 343634 31764 343640 31776
rect 343692 31764 343698 31816
rect 339736 31708 340920 31736
rect 339736 31696 339742 31708
rect 279418 31016 279424 31068
rect 279476 31056 279482 31068
rect 287698 31056 287704 31068
rect 279476 31028 287704 31056
rect 279476 31016 279482 31028
rect 287698 31016 287704 31028
rect 287756 31016 287762 31068
rect 338022 29792 338028 29844
rect 338080 29832 338086 29844
rect 339678 29832 339684 29844
rect 338080 29804 339684 29832
rect 338080 29792 338086 29804
rect 339678 29792 339684 29804
rect 339736 29792 339742 29844
rect 332594 27616 332600 27668
rect 332652 27656 332658 27668
rect 338022 27656 338028 27668
rect 332652 27628 338028 27656
rect 332652 27616 332658 27628
rect 338022 27616 338028 27628
rect 338080 27616 338086 27668
rect 551370 27548 551376 27600
rect 551428 27588 551434 27600
rect 580074 27588 580080 27600
rect 551428 27560 580080 27588
rect 551428 27548 551434 27560
rect 580074 27548 580080 27560
rect 580132 27548 580138 27600
rect 39574 25508 39580 25560
rect 39632 25548 39638 25560
rect 498194 25548 498200 25560
rect 39632 25520 498200 25548
rect 39632 25508 39638 25520
rect 498194 25508 498200 25520
rect 498252 25508 498258 25560
rect 331214 25304 331220 25356
rect 331272 25344 331278 25356
rect 335998 25344 336004 25356
rect 331272 25316 336004 25344
rect 331272 25304 331278 25316
rect 335998 25304 336004 25316
rect 336056 25304 336062 25356
rect 3234 24692 3240 24744
rect 3292 24732 3298 24744
rect 6362 24732 6368 24744
rect 3292 24704 6368 24732
rect 3292 24692 3298 24704
rect 6362 24692 6368 24704
rect 6420 24692 6426 24744
rect 326614 23536 326620 23588
rect 326672 23576 326678 23588
rect 331214 23576 331220 23588
rect 326672 23548 331220 23576
rect 326672 23536 326678 23548
rect 331214 23536 331220 23548
rect 331272 23536 331278 23588
rect 329834 23468 329840 23520
rect 329892 23508 329898 23520
rect 332594 23508 332600 23520
rect 329892 23480 332600 23508
rect 329892 23468 329898 23480
rect 332594 23468 332600 23480
rect 332652 23468 332658 23520
rect 326614 22148 326620 22160
rect 321572 22120 326620 22148
rect 320818 22040 320824 22092
rect 320876 22080 320882 22092
rect 321572 22080 321600 22120
rect 326614 22108 326620 22120
rect 326672 22108 326678 22160
rect 320876 22052 321600 22080
rect 320876 22040 320882 22052
rect 269114 19932 269120 19984
rect 269172 19972 269178 19984
rect 279418 19972 279424 19984
rect 269172 19944 279424 19972
rect 269172 19932 269178 19944
rect 279418 19932 279424 19944
rect 279476 19932 279482 19984
rect 61378 17892 61384 17944
rect 61436 17932 61442 17944
rect 64506 17932 64512 17944
rect 61436 17904 64512 17932
rect 61436 17892 61442 17904
rect 64506 17892 64512 17904
rect 64564 17892 64570 17944
rect 329466 15212 329472 15224
rect 327092 15184 329472 15212
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 11698 15144 11704 15156
rect 3476 15116 11704 15144
rect 3476 15104 3482 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 326338 15104 326344 15156
rect 326396 15144 326402 15156
rect 327092 15144 327120 15184
rect 329466 15172 329472 15184
rect 329524 15172 329530 15224
rect 340138 15172 340144 15224
rect 340196 15212 340202 15224
rect 341518 15212 341524 15224
rect 340196 15184 341524 15212
rect 340196 15172 340202 15184
rect 341518 15172 341524 15184
rect 341576 15172 341582 15224
rect 326396 15116 327120 15144
rect 326396 15104 326402 15116
rect 64506 10276 64512 10328
rect 64564 10316 64570 10328
rect 69658 10316 69664 10328
rect 64564 10288 69664 10316
rect 64564 10276 64570 10288
rect 69658 10276 69664 10288
rect 69716 10276 69722 10328
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 6270 9908 6276 9920
rect 3016 9880 6276 9908
rect 3016 9868 3022 9880
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 266170 8236 266176 8288
rect 266228 8276 266234 8288
rect 580166 8276 580172 8288
rect 266228 8248 580172 8276
rect 266228 8236 266234 8248
rect 580166 8236 580172 8248
rect 580224 8236 580230 8288
rect 376110 6264 376116 6316
rect 376168 6304 376174 6316
rect 545114 6304 545120 6316
rect 376168 6276 545120 6304
rect 376168 6264 376174 6276
rect 545114 6264 545120 6276
rect 545172 6264 545178 6316
rect 136358 6196 136364 6248
rect 136416 6236 136422 6248
rect 456794 6236 456800 6248
rect 136416 6208 456800 6236
rect 136416 6196 136422 6208
rect 456794 6196 456800 6208
rect 456852 6196 456858 6248
rect 93118 6128 93124 6180
rect 93176 6168 93182 6180
rect 542078 6168 542084 6180
rect 93176 6140 542084 6168
rect 93176 6128 93182 6140
rect 542078 6128 542084 6140
rect 542136 6128 542142 6180
rect 57882 5448 57888 5500
rect 57940 5488 57946 5500
rect 242894 5488 242900 5500
rect 57940 5460 242900 5488
rect 57940 5448 57946 5460
rect 242894 5448 242900 5460
rect 242952 5448 242958 5500
rect 282822 5448 282828 5500
rect 282880 5488 282886 5500
rect 544010 5488 544016 5500
rect 282880 5460 544016 5488
rect 282880 5448 282886 5460
rect 544010 5448 544016 5460
rect 544068 5448 544074 5500
rect 39850 5380 39856 5432
rect 39908 5420 39914 5432
rect 352742 5420 352748 5432
rect 39908 5392 352748 5420
rect 39908 5380 39914 5392
rect 352742 5380 352748 5392
rect 352800 5380 352806 5432
rect 356054 5380 356060 5432
rect 356112 5420 356118 5432
rect 545666 5420 545672 5432
rect 356112 5392 545672 5420
rect 356112 5380 356118 5392
rect 545666 5380 545672 5392
rect 545724 5380 545730 5432
rect 69750 5312 69756 5364
rect 69808 5352 69814 5364
rect 186314 5352 186320 5364
rect 69808 5324 186320 5352
rect 69808 5312 69814 5324
rect 186314 5312 186320 5324
rect 186372 5312 186378 5364
rect 229646 5312 229652 5364
rect 229704 5352 229710 5364
rect 542906 5352 542912 5364
rect 229704 5324 542912 5352
rect 229704 5312 229710 5324
rect 542906 5312 542912 5324
rect 542964 5312 542970 5364
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 4798 5284 4804 5296
rect 2832 5256 4804 5284
rect 2832 5244 2838 5256
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 79870 5244 79876 5296
rect 79928 5284 79934 5296
rect 396074 5284 396080 5296
rect 79928 5256 396080 5284
rect 79928 5244 79934 5256
rect 396074 5244 396080 5256
rect 396132 5244 396138 5296
rect 406102 5244 406108 5296
rect 406160 5284 406166 5296
rect 545482 5284 545488 5296
rect 406160 5256 545488 5284
rect 406160 5244 406166 5256
rect 545482 5244 545488 5256
rect 545540 5244 545546 5296
rect 37918 5176 37924 5228
rect 37976 5216 37982 5228
rect 409414 5216 409420 5228
rect 37976 5188 409420 5216
rect 37976 5176 37982 5188
rect 409414 5176 409420 5188
rect 409472 5176 409478 5228
rect 142982 5108 142988 5160
rect 143040 5148 143046 5160
rect 544102 5148 544108 5160
rect 143040 5120 544108 5148
rect 143040 5108 143046 5120
rect 544102 5108 544108 5120
rect 544160 5108 544166 5160
rect 39390 5040 39396 5092
rect 39448 5080 39454 5092
rect 452654 5080 452660 5092
rect 39448 5052 452660 5080
rect 39448 5040 39454 5052
rect 452654 5040 452660 5052
rect 452712 5040 452718 5092
rect 69658 4972 69664 5024
rect 69716 5012 69722 5024
rect 126422 5012 126428 5024
rect 69716 4984 126428 5012
rect 69716 4972 69722 4984
rect 126422 4972 126428 4984
rect 126480 4972 126486 5024
rect 129734 4972 129740 5024
rect 129792 5012 129798 5024
rect 545574 5012 545580 5024
rect 129792 4984 545580 5012
rect 129792 4972 129798 4984
rect 545574 4972 545580 4984
rect 545632 4972 545638 5024
rect 26510 4904 26516 4956
rect 26568 4944 26574 4956
rect 480254 4944 480260 4956
rect 26568 4916 480260 4944
rect 26568 4904 26574 4916
rect 480254 4904 480260 4916
rect 480312 4904 480318 4956
rect 49878 4836 49884 4888
rect 49936 4876 49942 4888
rect 541986 4876 541992 4888
rect 49936 4848 541992 4876
rect 49936 4836 49942 4848
rect 541986 4836 541992 4848
rect 542044 4836 542050 4888
rect 37458 4768 37464 4820
rect 37516 4808 37522 4820
rect 542446 4808 542452 4820
rect 37516 4780 542452 4808
rect 37516 4768 37522 4780
rect 542446 4768 542452 4780
rect 542504 4768 542510 4820
rect 111702 4700 111708 4752
rect 111760 4740 111766 4752
rect 256326 4740 256332 4752
rect 111760 4712 256332 4740
rect 111760 4700 111766 4712
rect 256326 4700 256332 4712
rect 256384 4700 256390 4752
rect 296254 4700 296260 4752
rect 296312 4740 296318 4752
rect 340138 4740 340144 4752
rect 296312 4712 340144 4740
rect 296312 4700 296318 4712
rect 340138 4700 340144 4712
rect 340196 4700 340202 4752
rect 389358 4700 389364 4752
rect 389416 4740 389422 4752
rect 505094 4740 505100 4752
rect 389416 4712 505100 4740
rect 389416 4700 389422 4712
rect 505094 4700 505100 4712
rect 505152 4700 505158 4752
rect 131022 4632 131028 4684
rect 131080 4672 131086 4684
rect 219710 4672 219716 4684
rect 131080 4644 219716 4672
rect 131080 4632 131086 4644
rect 219710 4632 219716 4644
rect 219768 4632 219774 4684
rect 226334 4632 226340 4684
rect 226392 4672 226398 4684
rect 299474 4672 299480 4684
rect 226392 4644 299480 4672
rect 226392 4632 226398 4644
rect 299474 4632 299480 4644
rect 299532 4632 299538 4684
rect 299566 4632 299572 4684
rect 299624 4672 299630 4684
rect 320818 4672 320824 4684
rect 299624 4644 320824 4672
rect 299624 4632 299630 4644
rect 320818 4632 320824 4644
rect 320876 4632 320882 4684
rect 357342 4632 357348 4684
rect 357400 4672 357406 4684
rect 442718 4672 442724 4684
rect 357400 4644 442724 4672
rect 357400 4632 357406 4644
rect 442718 4632 442724 4644
rect 442776 4632 442782 4684
rect 284294 4564 284300 4616
rect 284352 4604 284358 4616
rect 326338 4604 326344 4616
rect 284352 4576 326344 4604
rect 284352 4564 284358 4576
rect 326338 4564 326344 4576
rect 326396 4564 326402 4616
rect 41046 4088 41052 4140
rect 41104 4128 41110 4140
rect 183094 4128 183100 4140
rect 41104 4100 183100 4128
rect 41104 4088 41110 4100
rect 183094 4088 183100 4100
rect 183152 4088 183158 4140
rect 262950 4088 262956 4140
rect 263008 4128 263014 4140
rect 487154 4128 487160 4140
rect 263008 4100 487160 4128
rect 263008 4088 263014 4100
rect 487154 4088 487160 4100
rect 487212 4088 487218 4140
rect 539502 4088 539508 4140
rect 539560 4128 539566 4140
rect 575750 4128 575756 4140
rect 539560 4100 575756 4128
rect 539560 4088 539566 4100
rect 575750 4088 575756 4100
rect 575808 4088 575814 4140
rect 40678 4020 40684 4072
rect 40736 4060 40742 4072
rect 189718 4060 189724 4072
rect 40736 4032 189724 4060
rect 40736 4020 40742 4032
rect 189718 4020 189724 4032
rect 189776 4020 189782 4072
rect 206278 4020 206284 4072
rect 206336 4060 206342 4072
rect 219434 4060 219440 4072
rect 206336 4032 219440 4060
rect 206336 4020 206342 4032
rect 219434 4020 219440 4032
rect 219492 4020 219498 4072
rect 223022 4020 223028 4072
rect 223080 4060 223086 4072
rect 234614 4060 234620 4072
rect 223080 4032 234620 4060
rect 223080 4020 223086 4032
rect 234614 4020 234620 4032
rect 234672 4020 234678 4072
rect 255222 4020 255228 4072
rect 255280 4060 255286 4072
rect 492582 4060 492588 4072
rect 255280 4032 492588 4060
rect 255280 4020 255286 4032
rect 492582 4020 492588 4032
rect 492640 4020 492646 4072
rect 532602 4020 532608 4072
rect 532660 4060 532666 4072
rect 536837 4063 536895 4069
rect 536837 4060 536849 4063
rect 532660 4032 536849 4060
rect 532660 4020 532666 4032
rect 536837 4029 536849 4032
rect 536883 4029 536895 4063
rect 536837 4023 536895 4029
rect 542262 4020 542268 4072
rect 542320 4060 542326 4072
rect 579062 4060 579068 4072
rect 542320 4032 579068 4060
rect 542320 4020 542326 4032
rect 579062 4020 579068 4032
rect 579120 4020 579126 4072
rect 40218 3952 40224 4004
rect 40276 3992 40282 4004
rect 236270 3992 236276 4004
rect 40276 3964 236276 3992
rect 40276 3952 40282 3964
rect 236270 3952 236276 3964
rect 236328 3952 236334 4004
rect 276198 3952 276204 4004
rect 276256 3992 276262 4004
rect 277302 3992 277308 4004
rect 276256 3964 277308 3992
rect 276256 3952 276262 3964
rect 277302 3952 277308 3964
rect 277360 3952 277366 4004
rect 286134 3952 286140 4004
rect 286192 3992 286198 4004
rect 542538 3992 542544 4004
rect 286192 3964 542544 3992
rect 286192 3952 286198 3964
rect 542538 3952 542544 3964
rect 542596 3952 542602 4004
rect 547414 3952 547420 4004
rect 547472 3992 547478 4004
rect 580166 3992 580172 4004
rect 547472 3964 580172 3992
rect 547472 3952 547478 3964
rect 580166 3952 580172 3964
rect 580224 3952 580230 4004
rect 38562 3884 38568 3936
rect 38620 3924 38626 3936
rect 252830 3924 252836 3936
rect 38620 3896 252836 3924
rect 38620 3884 38626 3896
rect 252830 3884 252836 3896
rect 252888 3884 252894 3936
rect 272886 3884 272892 3936
rect 272944 3924 272950 3936
rect 277394 3924 277400 3936
rect 272944 3896 277400 3924
rect 272944 3884 272950 3896
rect 277394 3884 277400 3896
rect 277452 3884 277458 3936
rect 279510 3884 279516 3936
rect 279568 3924 279574 3936
rect 543090 3924 543096 3936
rect 279568 3896 543096 3924
rect 279568 3884 279574 3896
rect 543090 3884 543096 3896
rect 543148 3884 543154 3936
rect 40770 3816 40776 3868
rect 40828 3856 40834 3868
rect 319438 3856 319444 3868
rect 40828 3828 319444 3856
rect 40828 3816 40834 3828
rect 319438 3816 319444 3828
rect 319496 3816 319502 3868
rect 324222 3816 324228 3868
rect 324280 3856 324286 3868
rect 326062 3856 326068 3868
rect 324280 3828 326068 3856
rect 324280 3816 324286 3828
rect 326062 3816 326068 3828
rect 326120 3816 326126 3868
rect 400122 3816 400128 3868
rect 400180 3856 400186 3868
rect 582374 3856 582380 3868
rect 400180 3828 582380 3856
rect 400180 3816 400186 3828
rect 582374 3816 582380 3828
rect 582432 3816 582438 3868
rect 38010 3748 38016 3800
rect 38068 3788 38074 3800
rect 46566 3788 46572 3800
rect 38068 3760 46572 3788
rect 38068 3748 38074 3760
rect 46566 3748 46572 3760
rect 46624 3748 46630 3800
rect 59814 3748 59820 3800
rect 59872 3788 59878 3800
rect 340874 3788 340880 3800
rect 59872 3760 340880 3788
rect 59872 3748 59878 3760
rect 340874 3748 340880 3760
rect 340932 3748 340938 3800
rect 367738 3748 367744 3800
rect 367796 3788 367802 3800
rect 559190 3788 559196 3800
rect 367796 3760 559196 3788
rect 367796 3748 367802 3760
rect 559190 3748 559196 3760
rect 559248 3748 559254 3800
rect 39114 3680 39120 3732
rect 39172 3720 39178 3732
rect 322750 3720 322756 3732
rect 39172 3692 322756 3720
rect 39172 3680 39178 3692
rect 322750 3680 322756 3692
rect 322808 3680 322814 3732
rect 326982 3680 326988 3732
rect 327040 3720 327046 3732
rect 329558 3720 329564 3732
rect 327040 3692 329564 3720
rect 327040 3680 327046 3692
rect 329558 3680 329564 3692
rect 329616 3680 329622 3732
rect 332870 3680 332876 3732
rect 332928 3720 332934 3732
rect 333882 3720 333888 3732
rect 332928 3692 333888 3720
rect 332928 3680 332934 3692
rect 333882 3680 333888 3692
rect 333940 3680 333946 3732
rect 336182 3680 336188 3732
rect 336240 3720 336246 3732
rect 543182 3720 543188 3732
rect 336240 3692 543188 3720
rect 336240 3680 336246 3692
rect 543182 3680 543188 3692
rect 543240 3680 543246 3732
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 99374 3652 99380 3664
rect 3384 3624 99380 3652
rect 3384 3612 3390 3624
rect 99374 3612 99380 3624
rect 99432 3612 99438 3664
rect 113174 3612 113180 3664
rect 113232 3652 113238 3664
rect 140774 3652 140780 3664
rect 113232 3624 140780 3652
rect 113232 3612 113238 3624
rect 140774 3612 140780 3624
rect 140832 3612 140838 3664
rect 146478 3612 146484 3664
rect 146536 3652 146542 3664
rect 477494 3652 477500 3664
rect 146536 3624 477500 3652
rect 146536 3612 146542 3624
rect 477494 3612 477500 3624
rect 477552 3612 477558 3664
rect 505830 3612 505836 3664
rect 505888 3652 505894 3664
rect 542630 3652 542636 3664
rect 505888 3624 542636 3652
rect 505888 3612 505894 3624
rect 542630 3612 542636 3624
rect 542688 3612 542694 3664
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 153102 3584 153108 3596
rect 41288 3556 153108 3584
rect 41288 3544 41294 3556
rect 153102 3544 153108 3556
rect 153160 3544 153166 3596
rect 156414 3544 156420 3596
rect 156472 3584 156478 3596
rect 543550 3584 543556 3596
rect 156472 3556 543556 3584
rect 156472 3544 156478 3556
rect 543550 3544 543556 3556
rect 543608 3544 543614 3596
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13722 3516 13728 3528
rect 13320 3488 13728 3516
rect 13320 3476 13326 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17862 3516 17868 3528
rect 16632 3488 17868 3516
rect 16632 3476 16638 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 20622 3516 20628 3528
rect 19944 3488 20628 3516
rect 19944 3476 19950 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 34422 3516 34428 3528
rect 33192 3488 34428 3516
rect 33192 3476 33198 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 37090 3516 37096 3528
rect 36688 3488 37096 3516
rect 36688 3476 36694 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 43254 3476 43260 3528
rect 43312 3516 43318 3528
rect 44082 3516 44088 3528
rect 43312 3488 44088 3516
rect 43312 3476 43318 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 469214 3516 469220 3528
rect 44192 3488 469220 3516
rect 40494 3408 40500 3460
rect 40552 3448 40558 3460
rect 44192 3448 44220 3488
rect 469214 3476 469220 3488
rect 469272 3476 469278 3528
rect 495894 3476 495900 3528
rect 495952 3516 495958 3528
rect 545390 3516 545396 3528
rect 495952 3488 545396 3516
rect 495952 3476 495958 3488
rect 545390 3476 545396 3488
rect 545448 3476 545454 3528
rect 551278 3476 551284 3528
rect 551336 3516 551342 3528
rect 552566 3516 552572 3528
rect 551336 3488 552572 3516
rect 551336 3476 551342 3488
rect 552566 3476 552572 3488
rect 552624 3476 552630 3528
rect 552658 3476 552664 3528
rect 552716 3516 552722 3528
rect 569126 3516 569132 3528
rect 552716 3488 569132 3516
rect 552716 3476 552722 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 40552 3420 44220 3448
rect 44269 3451 44327 3457
rect 40552 3408 40558 3420
rect 44269 3417 44281 3451
rect 44315 3448 44327 3451
rect 522574 3448 522580 3460
rect 44315 3420 522580 3448
rect 44315 3417 44327 3420
rect 44269 3411 44327 3417
rect 522574 3408 522580 3420
rect 522632 3408 522638 3460
rect 535822 3408 535828 3460
rect 535880 3448 535886 3460
rect 536742 3448 536748 3460
rect 535880 3420 536748 3448
rect 535880 3408 535886 3420
rect 536742 3408 536748 3420
rect 536800 3408 536806 3460
rect 536837 3451 536895 3457
rect 536837 3417 536849 3451
rect 536883 3448 536895 3451
rect 572438 3448 572444 3460
rect 536883 3420 572444 3448
rect 536883 3417 536895 3420
rect 536837 3411 536895 3417
rect 572438 3408 572444 3420
rect 572496 3408 572502 3460
rect 40954 3340 40960 3392
rect 41012 3380 41018 3392
rect 166350 3380 166356 3392
rect 41012 3352 166356 3380
rect 41012 3340 41018 3352
rect 166350 3340 166356 3352
rect 166408 3340 166414 3392
rect 179598 3340 179604 3392
rect 179656 3380 179662 3392
rect 198734 3380 198740 3392
rect 179656 3352 198740 3380
rect 179656 3340 179662 3352
rect 198734 3340 198740 3352
rect 198792 3340 198798 3392
rect 263502 3340 263508 3392
rect 263560 3380 263566 3392
rect 485958 3380 485964 3392
rect 263560 3352 485964 3380
rect 263560 3340 263566 3352
rect 485958 3340 485964 3352
rect 486016 3340 486022 3392
rect 527082 3340 527088 3392
rect 527140 3380 527146 3392
rect 562502 3380 562508 3392
rect 527140 3352 562508 3380
rect 527140 3340 527146 3352
rect 562502 3340 562508 3352
rect 562560 3340 562566 3392
rect 38470 3272 38476 3324
rect 38528 3312 38534 3324
rect 44269 3315 44327 3321
rect 44269 3312 44281 3315
rect 38528 3284 44281 3312
rect 38528 3272 38534 3284
rect 44269 3281 44281 3284
rect 44315 3281 44327 3315
rect 44269 3275 44327 3281
rect 44361 3315 44419 3321
rect 44361 3281 44373 3315
rect 44407 3312 44419 3315
rect 47121 3315 47179 3321
rect 44407 3284 47072 3312
rect 44407 3281 44419 3284
rect 44361 3275 44419 3281
rect 40402 3204 40408 3256
rect 40460 3244 40466 3256
rect 46937 3247 46995 3253
rect 46937 3244 46949 3247
rect 40460 3216 46949 3244
rect 40460 3204 40466 3216
rect 46937 3213 46949 3216
rect 46983 3213 46995 3247
rect 47044 3244 47072 3284
rect 47121 3281 47133 3315
rect 47167 3312 47179 3315
rect 159726 3312 159732 3324
rect 47167 3284 159732 3312
rect 47167 3281 47179 3284
rect 47121 3275 47179 3281
rect 159726 3272 159732 3284
rect 159784 3272 159790 3324
rect 289446 3312 289452 3324
rect 161446 3284 289452 3312
rect 149790 3244 149796 3256
rect 47044 3216 149796 3244
rect 46937 3207 46995 3213
rect 149790 3204 149796 3216
rect 149848 3204 149854 3256
rect 159358 3204 159364 3256
rect 159416 3244 159422 3256
rect 161446 3244 161474 3284
rect 289446 3272 289452 3284
rect 289504 3272 289510 3324
rect 292942 3272 292948 3324
rect 293000 3312 293006 3324
rect 295426 3312 295432 3324
rect 293000 3284 295432 3312
rect 293000 3272 293006 3284
rect 295426 3272 295432 3284
rect 295484 3272 295490 3324
rect 312814 3272 312820 3324
rect 312872 3312 312878 3324
rect 517514 3312 517520 3324
rect 312872 3284 517520 3312
rect 312872 3272 312878 3284
rect 517514 3272 517520 3284
rect 517572 3272 517578 3324
rect 525886 3272 525892 3324
rect 525944 3312 525950 3324
rect 542998 3312 543004 3324
rect 525944 3284 543004 3312
rect 525944 3272 525950 3284
rect 542998 3272 543004 3284
rect 543056 3272 543062 3324
rect 159416 3216 161474 3244
rect 159416 3204 159422 3216
rect 186406 3204 186412 3256
rect 186464 3244 186470 3256
rect 187602 3244 187608 3256
rect 186464 3216 187608 3244
rect 186464 3204 186470 3216
rect 187602 3204 187608 3216
rect 187660 3204 187666 3256
rect 342806 3244 342812 3256
rect 187804 3216 342812 3244
rect 14 3136 20 3188
rect 72 3176 78 3188
rect 1302 3176 1308 3188
rect 72 3148 1308 3176
rect 72 3136 78 3148
rect 1302 3136 1308 3148
rect 1360 3136 1366 3188
rect 40862 3136 40868 3188
rect 40920 3176 40926 3188
rect 133046 3176 133052 3188
rect 40920 3148 133052 3176
rect 40920 3136 40926 3148
rect 133046 3136 133052 3148
rect 133104 3136 133110 3188
rect 176286 3136 176292 3188
rect 176344 3176 176350 3188
rect 187697 3179 187755 3185
rect 187697 3176 187709 3179
rect 176344 3148 187709 3176
rect 176344 3136 176350 3148
rect 187697 3145 187709 3148
rect 187743 3145 187755 3179
rect 187697 3139 187755 3145
rect 41690 3068 41696 3120
rect 41748 3108 41754 3120
rect 103054 3108 103060 3120
rect 41748 3080 103060 3108
rect 41748 3068 41754 3080
rect 103054 3068 103060 3080
rect 103112 3068 103118 3120
rect 131758 3068 131764 3120
rect 131816 3108 131822 3120
rect 163038 3108 163044 3120
rect 131816 3080 163044 3108
rect 131816 3068 131822 3080
rect 163038 3068 163044 3080
rect 163096 3068 163102 3120
rect 182818 3068 182824 3120
rect 182876 3108 182882 3120
rect 187804 3108 187832 3216
rect 342806 3204 342812 3216
rect 342864 3204 342870 3256
rect 360102 3204 360108 3256
rect 360160 3244 360166 3256
rect 366174 3244 366180 3256
rect 360160 3216 366180 3244
rect 360160 3204 360166 3216
rect 366174 3204 366180 3216
rect 366232 3204 366238 3256
rect 402882 3204 402888 3256
rect 402940 3244 402946 3256
rect 465902 3244 465908 3256
rect 402940 3216 465908 3244
rect 402940 3204 402946 3216
rect 465902 3204 465908 3216
rect 465960 3204 465966 3256
rect 532510 3204 532516 3256
rect 532568 3244 532574 3256
rect 545206 3244 545212 3256
rect 532568 3216 545212 3244
rect 532568 3204 532574 3216
rect 545206 3204 545212 3216
rect 545264 3204 545270 3256
rect 187881 3179 187939 3185
rect 187881 3145 187893 3179
rect 187927 3176 187939 3179
rect 193214 3176 193220 3188
rect 187927 3148 193220 3176
rect 187927 3145 187939 3148
rect 187881 3139 187939 3145
rect 193214 3136 193220 3148
rect 193272 3136 193278 3188
rect 202782 3136 202788 3188
rect 202840 3176 202846 3188
rect 346118 3176 346124 3188
rect 202840 3148 346124 3176
rect 202840 3136 202846 3148
rect 346118 3136 346124 3148
rect 346176 3136 346182 3188
rect 415302 3136 415308 3188
rect 415360 3176 415366 3188
rect 429286 3176 429292 3188
rect 415360 3148 429292 3176
rect 415360 3136 415366 3148
rect 429286 3136 429292 3148
rect 429344 3136 429350 3188
rect 439498 3136 439504 3188
rect 439556 3176 439562 3188
rect 446030 3176 446036 3188
rect 439556 3148 446036 3176
rect 439556 3136 439562 3148
rect 446030 3136 446036 3148
rect 446088 3136 446094 3188
rect 449342 3136 449348 3188
rect 449400 3176 449406 3188
rect 449802 3176 449808 3188
rect 449400 3148 449808 3176
rect 449400 3136 449406 3148
rect 449802 3136 449808 3148
rect 449860 3136 449866 3188
rect 451918 3136 451924 3188
rect 451976 3176 451982 3188
rect 455966 3176 455972 3188
rect 451976 3148 455972 3176
rect 451976 3136 451982 3148
rect 455966 3136 455972 3148
rect 456024 3136 456030 3188
rect 462590 3136 462596 3188
rect 462648 3176 462654 3188
rect 523034 3176 523040 3188
rect 462648 3148 523040 3176
rect 462648 3136 462654 3148
rect 523034 3136 523040 3148
rect 523092 3136 523098 3188
rect 306190 3108 306196 3120
rect 182876 3080 187832 3108
rect 190426 3080 306196 3108
rect 182876 3068 182882 3080
rect 23198 3000 23204 3052
rect 23256 3040 23262 3052
rect 58989 3043 59047 3049
rect 58989 3040 59001 3043
rect 23256 3012 59001 3040
rect 23256 3000 23262 3012
rect 58989 3009 59001 3012
rect 59035 3009 59047 3043
rect 58989 3003 59047 3009
rect 59081 3043 59139 3049
rect 59081 3009 59093 3043
rect 59127 3040 59139 3043
rect 64874 3040 64880 3052
rect 59127 3012 64880 3040
rect 59127 3009 59139 3012
rect 59081 3003 59139 3009
rect 64874 3000 64880 3012
rect 64932 3000 64938 3052
rect 76558 3000 76564 3052
rect 76616 3040 76622 3052
rect 131850 3040 131856 3052
rect 76616 3012 131856 3040
rect 76616 3000 76622 3012
rect 131850 3000 131856 3012
rect 131908 3000 131914 3052
rect 184842 3000 184848 3052
rect 184900 3040 184906 3052
rect 190426 3040 190454 3080
rect 306190 3068 306196 3080
rect 306248 3068 306254 3120
rect 311802 3068 311808 3120
rect 311860 3108 311866 3120
rect 399294 3108 399300 3120
rect 311860 3080 399300 3108
rect 311860 3068 311866 3080
rect 399294 3068 399300 3080
rect 399352 3068 399358 3120
rect 443638 3068 443644 3120
rect 443696 3108 443702 3120
rect 502518 3108 502524 3120
rect 443696 3080 502524 3108
rect 443696 3068 443702 3080
rect 502518 3068 502524 3080
rect 502576 3068 502582 3120
rect 184900 3012 190454 3040
rect 184900 3000 184906 3012
rect 199654 3000 199660 3052
rect 199712 3040 199718 3052
rect 284294 3040 284300 3052
rect 199712 3012 284300 3040
rect 199712 3000 199718 3012
rect 284294 3000 284300 3012
rect 284352 3000 284358 3052
rect 301498 3000 301504 3052
rect 301556 3040 301562 3052
rect 416038 3040 416044 3052
rect 301556 3012 416044 3040
rect 301556 3000 301562 3012
rect 416038 3000 416044 3012
rect 416096 3000 416102 3052
rect 448422 3000 448428 3052
rect 448480 3040 448486 3052
rect 472526 3040 472532 3052
rect 448480 3012 472532 3040
rect 448480 3000 448486 3012
rect 472526 3000 472532 3012
rect 472584 3000 472590 3052
rect 512638 3000 512644 3052
rect 512696 3040 512702 3052
rect 513282 3040 513288 3052
rect 512696 3012 513288 3040
rect 512696 3000 512702 3012
rect 513282 3000 513288 3012
rect 513340 3000 513346 3052
rect 39942 2932 39948 2984
rect 40000 2972 40006 2984
rect 77294 2972 77300 2984
rect 40000 2944 77300 2972
rect 40000 2932 40006 2944
rect 77294 2932 77300 2944
rect 77352 2932 77358 2984
rect 89806 2932 89812 2984
rect 89864 2972 89870 2984
rect 120074 2972 120080 2984
rect 89864 2944 120080 2972
rect 89864 2932 89870 2944
rect 120074 2932 120080 2944
rect 120132 2932 120138 2984
rect 123110 2932 123116 2984
rect 123168 2972 123174 2984
rect 147674 2972 147680 2984
rect 123168 2944 147680 2972
rect 123168 2932 123174 2944
rect 147674 2932 147680 2944
rect 147732 2932 147738 2984
rect 213822 2932 213828 2984
rect 213880 2972 213886 2984
rect 216214 2972 216220 2984
rect 213880 2944 216220 2972
rect 213880 2932 213886 2944
rect 216214 2932 216220 2944
rect 216272 2932 216278 2984
rect 29822 2864 29828 2916
rect 29880 2904 29886 2916
rect 59081 2907 59139 2913
rect 59081 2904 59093 2907
rect 29880 2876 59093 2904
rect 29880 2864 29886 2876
rect 59081 2873 59093 2876
rect 59127 2873 59139 2907
rect 59081 2867 59139 2873
rect 59173 2907 59231 2913
rect 59173 2873 59185 2907
rect 59219 2904 59231 2907
rect 62114 2904 62120 2916
rect 59219 2876 62120 2904
rect 59219 2873 59231 2876
rect 59173 2867 59231 2873
rect 62114 2864 62120 2876
rect 62172 2864 62178 2916
rect 63126 2864 63132 2916
rect 63184 2904 63190 2916
rect 92566 2904 92572 2916
rect 63184 2876 92572 2904
rect 63184 2864 63190 2876
rect 92566 2864 92572 2876
rect 92624 2864 92630 2916
rect 38654 2796 38660 2848
rect 38712 2836 38718 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 38712 2808 44373 2836
rect 38712 2796 38718 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 53190 2796 53196 2848
rect 53248 2836 53254 2848
rect 86954 2836 86960 2848
rect 53248 2808 86960 2836
rect 53248 2796 53254 2808
rect 86954 2796 86960 2808
rect 87012 2796 87018 2848
<< via1 >>
rect 314660 702992 314712 703044
rect 315948 702992 316000 703044
rect 3424 702448 3476 702500
rect 7748 702448 7800 702500
rect 38660 700952 38712 701004
rect 73068 700952 73120 701004
rect 73160 700952 73212 701004
rect 575572 700952 575624 701004
rect 40040 700884 40092 700936
rect 239404 700884 239456 700936
rect 302700 700884 302752 700936
rect 543924 700884 543976 700936
rect 38016 700816 38068 700868
rect 276020 700816 276072 700868
rect 299388 700816 299440 700868
rect 541992 700816 542044 700868
rect 37096 700748 37148 700800
rect 312636 700748 312688 700800
rect 329380 700748 329432 700800
rect 543832 700748 543884 700800
rect 41880 700680 41932 700732
rect 56324 700680 56376 700732
rect 62948 700680 63000 700732
rect 352472 700680 352524 700732
rect 352748 700680 352800 700732
rect 385868 700680 385920 700732
rect 398748 700680 398800 700732
rect 415860 700680 415912 700732
rect 419172 700680 419224 700732
rect 542268 700680 542320 700732
rect 38108 700612 38160 700664
rect 336004 700612 336056 700664
rect 345940 700612 345992 700664
rect 543740 700612 543792 700664
rect 38844 700544 38896 700596
rect 362500 700544 362552 700596
rect 395804 700544 395856 700596
rect 543648 700544 543700 700596
rect 37464 700476 37516 700528
rect 149612 700476 149664 700528
rect 166172 700476 166224 700528
rect 542820 700476 542872 700528
rect 39948 700408 40000 700460
rect 422484 700408 422536 700460
rect 455788 700408 455840 700460
rect 542176 700408 542228 700460
rect 547420 700408 547472 700460
rect 555700 700408 555752 700460
rect 39672 700340 39724 700392
rect 432420 700340 432472 700392
rect 459468 700340 459520 700392
rect 578884 700340 578936 700392
rect 38292 700272 38344 700324
rect 495716 700272 495768 700324
rect 508964 700272 509016 700324
rect 544200 700272 544252 700324
rect 550180 700272 550232 700324
rect 562324 700272 562376 700324
rect 39488 700204 39540 700256
rect 216036 700204 216088 700256
rect 236092 700204 236144 700256
rect 242164 700204 242216 700256
rect 282644 700204 282696 700256
rect 491944 700204 491996 700256
rect 40408 700136 40460 700188
rect 189540 700136 189592 700188
rect 256148 700136 256200 700188
rect 324320 700136 324372 700188
rect 325608 700136 325660 700188
rect 462412 700136 462464 700188
rect 464988 700136 465040 700188
rect 535644 700136 535696 700188
rect 9772 700068 9824 700120
rect 10968 700068 11020 700120
rect 26332 700068 26384 700120
rect 27528 700068 27580 700120
rect 41604 700068 41656 700120
rect 146300 700068 146352 700120
rect 169484 700068 169536 700120
rect 175924 700068 175976 700120
rect 202788 700068 202840 700120
rect 326804 700068 326856 700120
rect 352656 700068 352708 700120
rect 382556 700068 382608 700120
rect 416044 700068 416096 700120
rect 429108 700068 429160 700120
rect 461584 700068 461636 700120
rect 479156 700068 479208 700120
rect 485780 700068 485832 700120
rect 542912 700068 542964 700120
rect 41236 700000 41288 700052
rect 139492 700000 139544 700052
rect 152924 700000 152976 700052
rect 264980 700000 265032 700052
rect 489184 700000 489236 700052
rect 499028 700000 499080 700052
rect 39212 699932 39264 699984
rect 38384 699864 38436 699916
rect 43076 699864 43128 699916
rect 54484 699932 54536 699984
rect 159548 699932 159600 699984
rect 425796 699932 425848 699984
rect 426348 699932 426400 699984
rect 132868 699864 132920 699916
rect 150348 699864 150400 699916
rect 206100 699864 206152 699916
rect 36452 699796 36504 699848
rect 37188 699796 37240 699848
rect 41052 699796 41104 699848
rect 106188 699796 106240 699848
rect 112996 699796 113048 699848
rect 129004 699796 129056 699848
rect 142804 699796 142856 699848
rect 152464 699796 152516 699848
rect 3148 699728 3200 699780
rect 6184 699728 6236 699780
rect 41328 699728 41380 699780
rect 19708 699660 19760 699712
rect 20628 699660 20680 699712
rect 41788 699660 41840 699712
rect 46388 699660 46440 699712
rect 53012 699660 53064 699712
rect 53656 699660 53708 699712
rect 66904 699660 66956 699712
rect 69572 699660 69624 699712
rect 70308 699660 70360 699712
rect 76380 699728 76432 699780
rect 77208 699728 77260 699780
rect 83004 699728 83056 699780
rect 86316 699728 86368 699780
rect 86868 699728 86920 699780
rect 102876 699728 102928 699780
rect 109684 699728 109736 699780
rect 180064 699728 180116 699780
rect 182916 699728 182968 699780
rect 99564 699660 99616 699712
rect 119620 699660 119672 699712
rect 122104 699660 122156 699712
rect 122932 699660 122984 699712
rect 124128 699660 124180 699712
rect 172796 699660 172848 699712
rect 173808 699660 173860 699712
rect 179420 699660 179472 699712
rect 180708 699660 180760 699712
rect 196164 699660 196216 699712
rect 197268 699660 197320 699712
rect 199476 699660 199528 699712
rect 200028 699660 200080 699712
rect 212724 699660 212776 699712
rect 213828 699660 213880 699712
rect 219532 699660 219584 699712
rect 220728 699660 220780 699712
rect 222844 699660 222896 699712
rect 223488 699660 223540 699712
rect 259460 699660 259512 699712
rect 260748 699660 260800 699712
rect 269396 699660 269448 699712
rect 270408 699660 270460 699712
rect 272708 699660 272760 699712
rect 273168 699660 273220 699712
rect 278780 699660 278832 699712
rect 279332 699660 279384 699712
rect 289268 699660 289320 699712
rect 289728 699660 289780 699712
rect 309324 699660 309376 699712
rect 310428 699660 310480 699712
rect 352564 699660 352616 699712
rect 353208 699660 353260 699712
rect 436744 699660 436796 699712
rect 439228 699660 439280 699712
rect 465724 699660 465776 699712
rect 466368 699660 466420 699712
rect 505652 699660 505704 699712
rect 506388 699660 506440 699712
rect 512644 699660 512696 699712
rect 515772 699660 515824 699712
rect 519084 699660 519136 699712
rect 520188 699660 520240 699712
rect 326804 699592 326856 699644
rect 334624 699592 334676 699644
rect 29644 698912 29696 698964
rect 60004 698912 60056 698964
rect 68560 698912 68612 698964
rect 129556 698912 129608 698964
rect 264980 698640 265032 698692
rect 267004 698640 267056 698692
rect 3240 698300 3292 698352
rect 509884 698300 509936 698352
rect 64144 697552 64196 697604
rect 68560 697552 68612 697604
rect 244924 697552 244976 697604
rect 262772 697552 262824 697604
rect 285956 697552 286008 697604
rect 294604 697552 294656 697604
rect 109776 696192 109828 696244
rect 135904 696192 135956 696244
rect 324320 696192 324372 696244
rect 331864 696192 331916 696244
rect 3148 692792 3200 692844
rect 10324 692792 10376 692844
rect 294604 692724 294656 692776
rect 298008 692724 298060 692776
rect 334624 692588 334676 692640
rect 336464 692588 336516 692640
rect 544844 691364 544896 691416
rect 580172 691364 580224 691416
rect 331864 690004 331916 690056
rect 333244 690004 333296 690056
rect 336464 689732 336516 689784
rect 338764 689732 338816 689784
rect 298008 688984 298060 689036
rect 305092 688984 305144 689036
rect 62764 687420 62816 687472
rect 64144 687420 64196 687472
rect 267004 686468 267056 686520
rect 273260 686468 273312 686520
rect 552756 685856 552808 685908
rect 579620 685856 579672 685908
rect 234528 685108 234580 685160
rect 244924 685108 244976 685160
rect 305092 685108 305144 685160
rect 310244 685108 310296 685160
rect 273260 684496 273312 684548
rect 278872 684428 278924 684480
rect 310244 682592 310296 682644
rect 318708 682592 318760 682644
rect 278872 681708 278924 681760
rect 280804 681708 280856 681760
rect 338764 681708 338816 681760
rect 340144 681708 340196 681760
rect 333244 680892 333296 680944
rect 333980 680892 334032 680944
rect 332508 680348 332560 680400
rect 580172 680348 580224 680400
rect 318708 679600 318760 679652
rect 331864 679600 331916 679652
rect 61292 678988 61344 679040
rect 62764 678988 62816 679040
rect 228364 678240 228416 678292
rect 234528 678240 234580 678292
rect 333980 676812 334032 676864
rect 341524 676812 341576 676864
rect 171876 676336 171928 676388
rect 175280 676336 175332 676388
rect 59728 675792 59780 675844
rect 61292 675792 61344 675844
rect 166264 673480 166316 673532
rect 171876 673480 171928 673532
rect 341524 672528 341576 672580
rect 346308 672528 346360 672580
rect 280804 672052 280856 672104
rect 282920 671984 282972 672036
rect 331864 671304 331916 671356
rect 343640 671304 343692 671356
rect 554044 670692 554096 670744
rect 580172 670692 580224 670744
rect 340144 669332 340196 669384
rect 346124 669196 346176 669248
rect 282920 668584 282972 668636
rect 284944 668584 284996 668636
rect 222108 668108 222160 668160
rect 228364 668108 228416 668160
rect 57796 666544 57848 666596
rect 59728 666544 59780 666596
rect 548524 666544 548576 666596
rect 579620 666544 579672 666596
rect 64880 666476 64932 666528
rect 66904 666476 66956 666528
rect 98184 666476 98236 666528
rect 252560 666476 252612 666528
rect 270408 666476 270460 666528
rect 388812 666476 388864 666528
rect 161848 666408 161900 666460
rect 325700 666408 325752 666460
rect 340512 666408 340564 666460
rect 352748 666408 352800 666460
rect 353208 666408 353260 666460
rect 428188 666408 428240 666460
rect 197268 666340 197320 666392
rect 407120 666340 407172 666392
rect 70952 666272 71004 666324
rect 292580 666272 292632 666324
rect 316224 666272 316276 666324
rect 441620 666272 441672 666324
rect 136548 666204 136600 666256
rect 358636 666204 358688 666256
rect 422208 666204 422260 666256
rect 436744 666204 436796 666256
rect 122104 666136 122156 666188
rect 146484 666136 146536 666188
rect 164792 666136 164844 666188
rect 481640 666136 481692 666188
rect 79968 666068 80020 666120
rect 431316 666068 431368 666120
rect 492220 666068 492272 666120
rect 512644 666068 512696 666120
rect 124128 666000 124180 666052
rect 510068 666000 510120 666052
rect 86040 665932 86092 665984
rect 95240 665932 95292 665984
rect 134432 665932 134484 665984
rect 531320 665932 531372 665984
rect 39580 665864 39632 665916
rect 519084 665864 519136 665916
rect 52736 665796 52788 665848
rect 552020 665796 552072 665848
rect 167920 665728 167972 665780
rect 318800 665728 318852 665780
rect 346400 665728 346452 665780
rect 349068 665728 349120 665780
rect 86868 665660 86920 665712
rect 207204 665660 207256 665712
rect 223488 665660 223540 665712
rect 246580 665660 246632 665712
rect 193128 665592 193180 665644
rect 231308 665592 231360 665644
rect 214656 665184 214708 665236
rect 222108 665184 222160 665236
rect 49792 665116 49844 665168
rect 54484 665116 54536 665168
rect 113272 665116 113324 665168
rect 539600 665116 539652 665168
rect 5172 665048 5224 665100
rect 101036 665048 101088 665100
rect 107200 665048 107252 665100
rect 551284 665048 551336 665100
rect 38568 664980 38620 665032
rect 46572 664980 46624 665032
rect 60004 664980 60056 665032
rect 104164 664980 104216 665032
rect 135904 664980 135956 665032
rect 140412 664980 140464 665032
rect 176936 664980 176988 665032
rect 180064 664980 180116 665032
rect 249708 664980 249760 665032
rect 252560 664980 252612 665032
rect 266268 664980 266320 665032
rect 276756 664980 276808 665032
rect 304080 664980 304132 665032
rect 305000 664980 305052 665032
rect 331312 664980 331364 665032
rect 332508 664980 332560 665032
rect 337384 664980 337436 665032
rect 342260 664980 342312 665032
rect 373816 664980 373868 665032
rect 389180 664980 389232 665032
rect 413192 664980 413244 665032
rect 416044 664980 416096 665032
rect 458640 664980 458692 665032
rect 459468 664980 459520 665032
rect 473728 664980 473780 665032
rect 489184 664980 489236 665032
rect 491944 664980 491996 665032
rect 500960 664980 501012 665032
rect 509884 664980 509936 665032
rect 516140 664980 516192 665032
rect 10600 664912 10652 664964
rect 61660 664912 61712 664964
rect 70308 664912 70360 664964
rect 219164 664912 219216 664964
rect 234528 664912 234580 664964
rect 352656 664912 352708 664964
rect 361672 664912 361724 664964
rect 368480 664912 368532 664964
rect 385960 664912 386012 664964
rect 401600 664912 401652 664964
rect 466368 664912 466420 664964
rect 531320 664912 531372 664964
rect 7932 664844 7984 664896
rect 79876 664844 79928 664896
rect 89628 664844 89680 664896
rect 270684 664844 270736 664896
rect 289728 664844 289780 664896
rect 470692 664844 470744 664896
rect 482928 664844 482980 664896
rect 553032 664844 553084 664896
rect 5080 664776 5132 664828
rect 83004 664776 83056 664828
rect 119344 664776 119396 664828
rect 314660 664776 314712 664828
rect 352564 664776 352616 664828
rect 443460 664776 443512 664828
rect 446496 664776 446548 664828
rect 542360 664776 542412 664828
rect 27528 664708 27580 664760
rect 225236 664708 225288 664760
rect 242164 664708 242216 664760
rect 258540 664708 258592 664760
rect 273168 664708 273220 664760
rect 282920 664708 282972 664760
rect 334440 664708 334492 664760
rect 521660 664708 521712 664760
rect 522304 664708 522356 664760
rect 547604 664708 547656 664760
rect 9588 664640 9640 664692
rect 89076 664640 89128 664692
rect 109684 664640 109736 664692
rect 125324 664640 125376 664692
rect 129004 664640 129056 664692
rect 137468 664640 137520 664692
rect 189080 664640 189132 664692
rect 458180 664640 458232 664692
rect 476856 664640 476908 664692
rect 548892 664640 548944 664692
rect 3424 664572 3476 664624
rect 143540 664572 143592 664624
rect 152464 664572 152516 664624
rect 170772 664572 170824 664624
rect 10876 664504 10928 664556
rect 173716 664504 173768 664556
rect 9312 664436 9364 664488
rect 182916 664572 182968 664624
rect 455512 664572 455564 664624
rect 461584 664572 461636 664624
rect 485872 664572 485924 664624
rect 551376 664572 551428 664624
rect 176016 664504 176068 664556
rect 185860 664504 185912 664556
rect 186228 664504 186280 664556
rect 198004 664504 198056 664556
rect 210240 664504 210292 664556
rect 558920 664504 558972 664556
rect 180708 664436 180760 664488
rect 534172 664436 534224 664488
rect 537392 664436 537444 664488
rect 545120 664436 545172 664488
rect 6552 664368 6604 664420
rect 195060 664368 195112 664420
rect 11704 664300 11756 664352
rect 249524 664300 249576 664352
rect 264704 664300 264756 664352
rect 336740 664368 336792 664420
rect 370688 664368 370740 664420
rect 375380 664368 375432 664420
rect 376760 664368 376812 664420
rect 391940 664368 391992 664420
rect 416136 664368 416188 664420
rect 549996 664368 550048 664420
rect 349528 664300 349580 664352
rect 548708 664300 548760 664352
rect 9404 664232 9456 664284
rect 267740 664232 267792 664284
rect 322296 664232 322348 664284
rect 551836 664232 551888 664284
rect 4988 664164 5040 664216
rect 288900 664164 288952 664216
rect 291936 664164 291988 664216
rect 551560 664164 551612 664216
rect 7656 664096 7708 664148
rect 313280 664096 313332 664148
rect 319352 664096 319404 664148
rect 549260 664096 549312 664148
rect 4804 664028 4856 664080
rect 222384 664028 222436 664080
rect 552848 664028 552900 664080
rect 10416 663960 10468 664012
rect 204076 663960 204128 664012
rect 213184 663960 213236 664012
rect 548800 663960 548852 664012
rect 3424 663892 3476 663944
rect 10508 663892 10560 663944
rect 10692 663892 10744 663944
rect 382740 663892 382792 663944
rect 548984 663892 549036 663944
rect 4712 663824 4764 663876
rect 131396 663824 131448 663876
rect 173808 663824 173860 663876
rect 38476 663756 38528 663808
rect 43628 663756 43680 663808
rect 142160 663756 142212 663808
rect 152556 663756 152608 663808
rect 228364 663756 228416 663808
rect 364800 663756 364852 663808
rect 494796 663824 494848 663876
rect 507032 663824 507084 663876
rect 550272 663824 550324 663876
rect 488816 663756 488868 663808
rect 491300 663756 491352 663808
rect 540336 663756 540388 663808
rect 542452 663756 542504 663808
rect 336740 663688 336792 663740
rect 353300 663688 353352 663740
rect 355968 663688 356020 663740
rect 546868 663688 546920 663740
rect 260748 663620 260800 663672
rect 542728 663620 542780 663672
rect 261760 663552 261812 663604
rect 580448 663552 580500 663604
rect 5264 663484 5316 663536
rect 328276 663484 328328 663536
rect 339408 663484 339460 663536
rect 543372 663484 543424 663536
rect 122472 663459 122524 663468
rect 122472 663425 122481 663459
rect 122481 663425 122515 663459
rect 122515 663425 122524 663459
rect 122472 663416 122524 663425
rect 213828 663416 213880 663468
rect 546684 663416 546736 663468
rect 39304 663348 39356 663400
rect 372620 663348 372672 663400
rect 59268 663280 59320 663332
rect 142160 663280 142212 663332
rect 209688 663280 209740 663332
rect 545396 663280 545448 663332
rect 41144 663212 41196 663264
rect 378140 663212 378192 663264
rect 40132 663144 40184 663196
rect 434720 663144 434772 663196
rect 77208 663076 77260 663128
rect 544016 663076 544068 663128
rect 53656 663008 53708 663060
rect 546500 663008 546552 663060
rect 9496 662940 9548 662992
rect 403716 662940 403768 662992
rect 5448 662872 5500 662924
rect 409880 662872 409932 662924
rect 5356 662804 5408 662856
rect 418804 662804 418856 662856
rect 433892 662847 433944 662856
rect 433892 662813 433901 662847
rect 433901 662813 433935 662847
rect 433935 662813 433944 662847
rect 433892 662804 433944 662813
rect 479340 662847 479392 662856
rect 479340 662813 479349 662847
rect 479349 662813 479383 662847
rect 479383 662813 479392 662847
rect 479340 662804 479392 662813
rect 95148 662736 95200 662788
rect 547144 662736 547196 662788
rect 77208 662711 77260 662720
rect 77208 662677 77217 662711
rect 77217 662677 77251 662711
rect 77251 662677 77260 662711
rect 77208 662668 77260 662677
rect 110420 662711 110472 662720
rect 110420 662677 110429 662711
rect 110429 662677 110463 662711
rect 110463 662677 110472 662711
rect 110420 662668 110472 662677
rect 116768 662668 116820 662720
rect 580356 662668 580408 662720
rect 49884 662643 49936 662652
rect 49884 662609 49893 662643
rect 49893 662609 49927 662643
rect 49927 662609 49936 662643
rect 49884 662600 49936 662609
rect 59912 662643 59964 662652
rect 59912 662609 59921 662643
rect 59921 662609 59955 662643
rect 59955 662609 59964 662643
rect 59912 662600 59964 662609
rect 68192 662600 68244 662652
rect 548616 662600 548668 662652
rect 9128 662532 9180 662584
rect 497556 662532 497608 662584
rect 506388 662575 506440 662584
rect 506388 662541 506397 662575
rect 506397 662541 506431 662575
rect 506431 662541 506440 662575
rect 506388 662532 506440 662541
rect 40592 662328 40644 662380
rect 543464 662464 543516 662516
rect 544108 662396 544160 662448
rect 125600 662328 125652 662380
rect 155960 662328 156012 662380
rect 354036 662371 354088 662380
rect 354036 662337 354045 662371
rect 354045 662337 354079 662371
rect 354079 662337 354088 662371
rect 354036 662328 354088 662337
rect 358268 662371 358320 662380
rect 358268 662337 358277 662371
rect 358277 662337 358311 662371
rect 358311 662337 358320 662371
rect 358268 662328 358320 662337
rect 425060 662371 425112 662380
rect 425060 662337 425069 662371
rect 425069 662337 425103 662371
rect 425103 662337 425112 662371
rect 425060 662328 425112 662337
rect 426348 662328 426400 662380
rect 546776 662328 546828 662380
rect 38936 662260 38988 662312
rect 241520 662260 241572 662312
rect 310428 662260 310480 662312
rect 545672 662260 545724 662312
rect 40684 662192 40736 662244
rect 158536 662192 158588 662244
rect 220728 662192 220780 662244
rect 542636 662192 542688 662244
rect 40500 662124 40552 662176
rect 245752 662124 245804 662176
rect 286416 662124 286468 662176
rect 545764 662124 545816 662176
rect 8116 662056 8168 662108
rect 128360 662056 128412 662108
rect 155868 662099 155920 662108
rect 155868 662065 155877 662099
rect 155877 662065 155911 662099
rect 155911 662065 155920 662099
rect 155868 662056 155920 662065
rect 200028 662056 200080 662108
rect 545488 662056 545540 662108
rect 7840 661988 7892 662040
rect 309692 661988 309744 662040
rect 346952 661988 347004 662040
rect 545212 661988 545264 662040
rect 6644 661920 6696 661972
rect 200764 661920 200816 661972
rect 216588 661920 216640 661972
rect 580264 661920 580316 661972
rect 37832 661852 37884 661904
rect 471980 661852 472032 661904
rect 476028 661852 476080 661904
rect 545948 661852 546000 661904
rect 4896 661784 4948 661836
rect 379520 661784 379572 661836
rect 392400 661784 392452 661836
rect 547328 661784 547380 661836
rect 4068 661716 4120 661768
rect 400588 661716 400640 661768
rect 412548 661716 412600 661768
rect 545580 661716 545632 661768
rect 37556 661648 37608 661700
rect 512000 661648 512052 661700
rect 515220 661691 515272 661700
rect 515220 661657 515229 661691
rect 515229 661657 515263 661691
rect 515263 661657 515272 661691
rect 515220 661648 515272 661657
rect 520188 661691 520240 661700
rect 520188 661657 520197 661691
rect 520197 661657 520231 661691
rect 520231 661657 520240 661691
rect 520188 661648 520240 661657
rect 539600 661648 539652 661700
rect 580724 661648 580776 661700
rect 3240 661580 3292 661632
rect 543280 661580 543332 661632
rect 6368 661512 6420 661564
rect 580540 661512 580592 661564
rect 3976 661444 4028 661496
rect 543096 661444 543148 661496
rect 40224 661376 40276 661428
rect 543004 661376 543056 661428
rect 37372 661240 37424 661292
rect 41696 661308 41748 661360
rect 542268 661308 542320 661360
rect 544384 661308 544436 661360
rect 35900 661172 35952 661224
rect 3608 661104 3660 661156
rect 544568 661240 544620 661292
rect 542084 661172 542136 661224
rect 544752 661104 544804 661156
rect 551468 661104 551520 661156
rect 579620 661104 579672 661156
rect 39856 661036 39908 661088
rect 565820 661036 565872 661088
rect 6828 660968 6880 661020
rect 38752 660968 38804 661020
rect 37924 660900 37976 660952
rect 41696 660968 41748 661020
rect 40316 660900 40368 660952
rect 37648 660832 37700 660884
rect 39304 660807 39356 660816
rect 39304 660773 39313 660807
rect 39313 660773 39347 660807
rect 39347 660773 39356 660807
rect 39304 660764 39356 660773
rect 41420 660764 41472 660816
rect 541900 660875 541952 660884
rect 541900 660841 541909 660875
rect 541909 660841 541943 660875
rect 541943 660841 541952 660875
rect 541900 660832 541952 660841
rect 542268 660764 542320 660816
rect 38200 660696 38252 660748
rect 541900 660696 541952 660748
rect 543556 660628 543608 660680
rect 39304 660560 39356 660612
rect 542544 660560 542596 660612
rect 40132 660492 40184 660544
rect 40776 660492 40828 660544
rect 545304 660492 545356 660544
rect 39028 660424 39080 660476
rect 568580 660424 568632 660476
rect 37004 660356 37056 660408
rect 40592 660356 40644 660408
rect 40868 660356 40920 660408
rect 580632 660356 580684 660408
rect 3884 660288 3936 660340
rect 544936 660288 544988 660340
rect 37280 660220 37332 660272
rect 542084 660220 542136 660272
rect 542544 660220 542596 660272
rect 542728 660220 542780 660272
rect 543464 660220 543516 660272
rect 39580 660152 39632 660204
rect 543188 660152 543240 660204
rect 39120 660084 39172 660136
rect 543464 660084 543516 660136
rect 544016 660084 544068 660136
rect 37740 660016 37792 660068
rect 545028 660016 545080 660068
rect 39764 659948 39816 660000
rect 549076 659948 549128 660000
rect 23480 659880 23532 659932
rect 544476 659880 544528 659932
rect 6460 659812 6512 659864
rect 544016 659812 544068 659864
rect 40132 659744 40184 659796
rect 580172 659744 580224 659796
rect 3332 659676 3384 659728
rect 546592 659676 546644 659728
rect 542728 659608 542780 659660
rect 543372 659608 543424 659660
rect 544660 659608 544712 659660
rect 581000 659608 581052 659660
rect 543372 659515 543424 659524
rect 543372 659481 543381 659515
rect 543381 659481 543415 659515
rect 543415 659481 543424 659515
rect 543372 659472 543424 659481
rect 544108 659268 544160 659320
rect 544752 659268 544804 659320
rect 544108 659175 544160 659184
rect 544108 659141 544117 659175
rect 544117 659141 544151 659175
rect 544151 659141 544160 659175
rect 544108 659132 544160 659141
rect 40592 658656 40644 658708
rect 41144 658656 41196 658708
rect 3424 658384 3476 658436
rect 6736 658384 6788 658436
rect 38844 658384 38896 658436
rect 32220 658180 32272 658232
rect 37004 658248 37056 658300
rect 34520 658180 34572 658232
rect 37740 658248 37792 658300
rect 37372 658112 37424 658164
rect 37740 658112 37792 658164
rect 38844 658044 38896 658096
rect 41144 657364 41196 657416
rect 41420 657364 41472 657416
rect 39304 657271 39356 657280
rect 39304 657237 39313 657271
rect 39313 657237 39347 657271
rect 39347 657237 39356 657271
rect 39304 657228 39356 657237
rect 41420 657271 41472 657280
rect 41420 657237 41429 657271
rect 41429 657237 41463 657271
rect 41463 657237 41472 657271
rect 41420 657228 41472 657237
rect 31024 657160 31076 657212
rect 35808 657160 35860 657212
rect 38936 657160 38988 657212
rect 40316 657160 40368 657212
rect 36912 657024 36964 657076
rect 37280 657024 37332 657076
rect 40316 657067 40368 657076
rect 40316 657033 40325 657067
rect 40325 657033 40359 657067
rect 40359 657033 40368 657067
rect 40316 657024 40368 657033
rect 19984 656888 20036 656940
rect 23480 656888 23532 656940
rect 544108 655596 544160 655648
rect 29828 655460 29880 655512
rect 32220 655528 32272 655580
rect 543648 655460 543700 655512
rect 544108 655460 544160 655512
rect 38844 655324 38896 655376
rect 40960 655324 41012 655376
rect 40776 655188 40828 655240
rect 40960 655188 41012 655240
rect 544016 655052 544068 655104
rect 544292 655052 544344 655104
rect 544292 654916 544344 654968
rect 544568 654916 544620 654968
rect 544568 654823 544620 654832
rect 544568 654789 544577 654823
rect 544577 654789 544611 654823
rect 544611 654789 544620 654823
rect 544568 654780 544620 654789
rect 33140 654576 33192 654628
rect 34520 654576 34572 654628
rect 3424 654440 3476 654492
rect 7564 654440 7616 654492
rect 3608 654372 3660 654424
rect 3424 654304 3476 654356
rect 542176 654347 542228 654356
rect 542176 654313 542185 654347
rect 542185 654313 542219 654347
rect 542219 654313 542228 654347
rect 542176 654304 542228 654313
rect 3240 654236 3292 654288
rect 3608 654236 3660 654288
rect 541900 654236 541952 654288
rect 32956 654168 33008 654220
rect 36912 654168 36964 654220
rect 40684 653964 40736 654016
rect 41420 654100 41472 654152
rect 541900 654143 541952 654146
rect 541900 654109 541909 654143
rect 541909 654109 541943 654143
rect 541943 654109 541952 654143
rect 541900 654094 541952 654109
rect 542084 654100 542136 654152
rect 37372 652740 37424 652792
rect 38844 652740 38896 652792
rect 40684 652740 40736 652792
rect 17960 651380 18012 651432
rect 19984 651380 20036 651432
rect 29000 651380 29052 651432
rect 31024 651380 31076 651432
rect 562324 651380 562376 651432
rect 3516 651312 3568 651364
rect 38844 651312 38896 651364
rect 567844 651312 567896 651364
rect 543648 651244 543700 651296
rect 38844 650700 38896 650752
rect 26700 650020 26752 650072
rect 29828 650020 29880 650072
rect 27068 648728 27120 648780
rect 29000 648728 29052 648780
rect 567844 648592 567896 648644
rect 36912 648524 36964 648576
rect 37372 648524 37424 648576
rect 571984 648524 572036 648576
rect 37280 648456 37332 648508
rect 38844 648456 38896 648508
rect 28264 647504 28316 647556
rect 33140 647504 33192 647556
rect 31484 647232 31536 647284
rect 32956 647232 33008 647284
rect 3700 647164 3752 647216
rect 38844 647164 38896 647216
rect 24952 645940 25004 645992
rect 27068 645940 27120 645992
rect 13820 645872 13872 645924
rect 17868 645872 17920 645924
rect 22100 645804 22152 645856
rect 26700 645872 26752 645924
rect 34520 645872 34572 645924
rect 36912 645872 36964 645924
rect 29920 645192 29972 645244
rect 31484 645192 31536 645244
rect 37372 643152 37424 643204
rect 38844 643152 38896 643204
rect 30380 643084 30432 643136
rect 34520 643084 34572 643136
rect 34612 643084 34664 643136
rect 37280 643084 37332 643136
rect 3792 643016 3844 643068
rect 38844 643016 38896 643068
rect 550088 641724 550140 641776
rect 580080 641724 580132 641776
rect 27620 640364 27672 640416
rect 30380 640364 30432 640416
rect 22744 640296 22796 640348
rect 24952 640296 25004 640348
rect 28172 640296 28224 640348
rect 29920 640296 29972 640348
rect 2780 640228 2832 640280
rect 4896 640228 4948 640280
rect 11060 638936 11112 638988
rect 13728 638936 13780 638988
rect 32956 638936 33008 638988
rect 34612 638936 34664 638988
rect 8484 637508 8536 637560
rect 11060 637576 11112 637628
rect 544844 637508 544896 637560
rect 580908 637508 580960 637560
rect 20260 637304 20312 637356
rect 22008 637304 22060 637356
rect 26240 637304 26292 637356
rect 28172 637304 28224 637356
rect 35256 636148 35308 636200
rect 37924 636216 37976 636268
rect 563704 636216 563756 636268
rect 579988 636216 580040 636268
rect 30380 635128 30432 635180
rect 32956 635128 33008 635180
rect 5540 634720 5592 634772
rect 8484 634788 8536 634840
rect 23480 634720 23532 634772
rect 27528 634788 27580 634840
rect 2780 633496 2832 633548
rect 4896 633496 4948 633548
rect 30104 633360 30156 633412
rect 35164 633428 35216 633480
rect 17224 632068 17276 632120
rect 20260 632068 20312 632120
rect 19156 632000 19208 632052
rect 23480 632068 23532 632120
rect 24860 631320 24912 631372
rect 30288 631320 30340 631372
rect 3516 630572 3568 630624
rect 7656 630572 7708 630624
rect 21364 630572 21416 630624
rect 26148 630640 26200 630692
rect 26884 630640 26936 630692
rect 30104 630640 30156 630692
rect 544108 629960 544160 630012
rect 544844 629960 544896 630012
rect 4620 629892 4672 629944
rect 5540 629892 5592 629944
rect 15844 629620 15896 629672
rect 19156 629620 19208 629672
rect 571984 629212 572036 629264
rect 575480 629212 575532 629264
rect 22100 627376 22152 627428
rect 24768 627376 24820 627428
rect 575480 626560 575532 626612
rect 576860 626560 576912 626612
rect 33784 626492 33836 626544
rect 35256 626492 35308 626544
rect 32404 625200 32456 625252
rect 37372 625200 37424 625252
rect 17960 623840 18012 623892
rect 22744 623840 22796 623892
rect 19984 623772 20036 623824
rect 22100 623772 22152 623824
rect 549076 623704 549128 623756
rect 580172 623704 580224 623756
rect 8208 622344 8260 622396
rect 15844 622412 15896 622464
rect 576860 621460 576912 621512
rect 579528 621460 579580 621512
rect 20076 620984 20128 621036
rect 21364 620984 21416 621036
rect 542268 620304 542320 620356
rect 542636 620304 542688 620356
rect 15844 619556 15896 619608
rect 17224 619556 17276 619608
rect 21364 619556 21416 619608
rect 26884 619556 26936 619608
rect 3792 619488 3844 619540
rect 8208 619488 8260 619540
rect 14464 619488 14516 619540
rect 17868 619488 17920 619540
rect 25504 618264 25556 618316
rect 38844 618264 38896 618316
rect 544844 618264 544896 618316
rect 578884 618264 578936 618316
rect 3516 618196 3568 618248
rect 4620 618196 4672 618248
rect 549904 616836 549956 616888
rect 579988 616836 580040 616888
rect 3332 615408 3384 615460
rect 32404 615408 32456 615460
rect 13820 614116 13872 614168
rect 15844 614116 15896 614168
rect 18052 614116 18104 614168
rect 20076 614116 20128 614168
rect 18788 614048 18840 614100
rect 21364 614116 21416 614168
rect 22100 614116 22152 614168
rect 28264 614116 28316 614168
rect 29644 614116 29696 614168
rect 38844 614116 38896 614168
rect 546960 613368 547012 613420
rect 580816 613368 580868 613420
rect 15844 611124 15896 611176
rect 18052 611124 18104 611176
rect 3332 610104 3384 610156
rect 8852 610104 8904 610156
rect 9036 609900 9088 609952
rect 18788 609968 18840 610020
rect 11336 608200 11388 608252
rect 13728 608200 13780 608252
rect 550364 607180 550416 607232
rect 580172 607180 580224 607232
rect 17960 607112 18012 607164
rect 19984 607112 20036 607164
rect 20168 606704 20220 606756
rect 22008 606704 22060 606756
rect 544844 605956 544896 606008
rect 546960 605956 547012 606008
rect 15200 605072 15252 605124
rect 20168 605072 20220 605124
rect 13820 604596 13872 604648
rect 17960 604596 18012 604648
rect 8208 604528 8260 604580
rect 11336 604528 11388 604580
rect 13912 604528 13964 604580
rect 15844 604528 15896 604580
rect 3332 604460 3384 604512
rect 21364 604460 21416 604512
rect 548984 604392 549036 604444
rect 579620 604392 579672 604444
rect 29736 603100 29788 603152
rect 33784 603100 33836 603152
rect 11428 601740 11480 601792
rect 13912 601740 13964 601792
rect 10968 601672 11020 601724
rect 13820 601672 13872 601724
rect 3700 601604 3752 601656
rect 38844 601604 38896 601656
rect 2780 601332 2832 601384
rect 4712 601332 4764 601384
rect 543556 600924 543608 600976
rect 558276 600924 558328 600976
rect 7656 600244 7708 600296
rect 9036 600244 9088 600296
rect 13084 600244 13136 600296
rect 15200 600312 15252 600364
rect 5540 597524 5592 597576
rect 8208 597524 8260 597576
rect 558184 597524 558236 597576
rect 580172 597524 580224 597576
rect 6736 597456 6788 597508
rect 38844 597456 38896 597508
rect 558276 597456 558328 597508
rect 562968 597456 563020 597508
rect 543648 596980 543700 597032
rect 550088 596980 550140 597032
rect 10784 596776 10836 596828
rect 11428 596776 11480 596828
rect 3332 595008 3384 595060
rect 9220 595008 9272 595060
rect 10232 594804 10284 594856
rect 13084 594804 13136 594856
rect 3332 593376 3384 593428
rect 5540 593376 5592 593428
rect 562968 593308 563020 593360
rect 579620 593308 579672 593360
rect 33784 592016 33836 592068
rect 38844 592016 38896 592068
rect 8300 591064 8352 591116
rect 10232 591064 10284 591116
rect 8024 590588 8076 590640
rect 10968 590656 11020 590708
rect 3148 590316 3200 590368
rect 6552 590316 6604 590368
rect 3884 589228 3936 589280
rect 38844 589228 38896 589280
rect 28264 587936 28316 587988
rect 29736 587936 29788 587988
rect 548984 587868 549036 587920
rect 580172 587868 580224 587920
rect 9680 586440 9732 586492
rect 14464 586508 14516 586560
rect 2780 585760 2832 585812
rect 4988 585760 5040 585812
rect 3240 585148 3292 585200
rect 8208 585148 8260 585200
rect 9036 583720 9088 583772
rect 9680 583720 9732 583772
rect 38936 582836 38988 582888
rect 40684 582836 40736 582888
rect 4160 582292 4212 582344
rect 8024 582360 8076 582412
rect 545856 582360 545908 582412
rect 579988 582360 580040 582412
rect 4252 580932 4304 580984
rect 7656 581000 7708 581052
rect 3700 579640 3752 579692
rect 4160 579640 4212 579692
rect 548892 579572 548944 579624
rect 579620 579572 579672 579624
rect 3240 578688 3292 578740
rect 4252 578688 4304 578740
rect 545304 578212 545356 578264
rect 567844 578212 567896 578264
rect 8300 577124 8352 577176
rect 10784 577124 10836 577176
rect 26884 575492 26936 575544
rect 28264 575492 28316 575544
rect 545028 574880 545080 574932
rect 544936 574676 544988 574728
rect 550364 574676 550416 574728
rect 544936 574540 544988 574592
rect 8024 574132 8076 574184
rect 9036 574132 9088 574184
rect 4988 574064 5040 574116
rect 38844 574064 38896 574116
rect 4712 573724 4764 573776
rect 8300 573724 8352 573776
rect 547236 572704 547288 572756
rect 580172 572704 580224 572756
rect 3056 570256 3108 570308
rect 7656 570256 7708 570308
rect 39120 568964 39172 569016
rect 41512 568964 41564 569016
rect 4344 568488 4396 568540
rect 8024 568556 8076 568608
rect 25596 568556 25648 568608
rect 26884 568556 26936 568608
rect 2780 565972 2832 566024
rect 5448 565972 5500 566024
rect 3056 565836 3108 565888
rect 4344 565836 4396 565888
rect 544936 565768 544988 565820
rect 580632 565768 580684 565820
rect 3884 564408 3936 564460
rect 4712 564408 4764 564460
rect 39948 562300 40000 562352
rect 40224 562300 40276 562352
rect 3148 561620 3200 561672
rect 38660 561620 38712 561672
rect 3148 560260 3200 560312
rect 14464 560260 14516 560312
rect 21732 559784 21784 559836
rect 25596 559784 25648 559836
rect 548708 558832 548760 558884
rect 580172 558832 580224 558884
rect 24124 556180 24176 556232
rect 38660 556180 38712 556232
rect 3148 556112 3200 556164
rect 21732 556112 21784 556164
rect 556804 553392 556856 553444
rect 580172 553392 580224 553444
rect 544936 552100 544988 552152
rect 548984 552100 549036 552152
rect 3148 550740 3200 550792
rect 6552 550740 6604 550792
rect 39948 548972 40000 549024
rect 41328 548972 41380 549024
rect 544660 547680 544712 547732
rect 544936 547680 544988 547732
rect 543464 547136 543516 547188
rect 546040 547136 546092 547188
rect 544660 546456 544712 546508
rect 562324 546456 562376 546508
rect 542176 543192 542228 543244
rect 543464 543192 543516 543244
rect 3148 540948 3200 541000
rect 35164 540948 35216 541000
rect 7748 539520 7800 539572
rect 38660 539520 38712 539572
rect 548708 538840 548760 538892
rect 580080 538840 580132 538892
rect 559564 538228 559616 538280
rect 580172 538228 580224 538280
rect 546040 537480 546092 537532
rect 553400 537480 553452 537532
rect 544660 535372 544712 535424
rect 554044 535372 554096 535424
rect 553400 533332 553452 533384
rect 565084 533332 565136 533384
rect 2780 531224 2832 531276
rect 5356 531224 5408 531276
rect 6736 529932 6788 529984
rect 38660 529932 38712 529984
rect 550456 528572 550508 528624
rect 580172 528572 580224 528624
rect 565084 527076 565136 527128
rect 569040 527076 569092 527128
rect 21364 525716 21416 525768
rect 38660 525716 38712 525768
rect 569040 522928 569092 522980
rect 571984 522928 572036 522980
rect 577504 521160 577556 521212
rect 579620 521160 579672 521212
rect 544660 520820 544712 520872
rect 548708 520820 548760 520872
rect 3148 520276 3200 520328
rect 21364 520276 21416 520328
rect 571984 518168 572036 518220
rect 580172 518168 580224 518220
rect 3148 516672 3200 516724
rect 3700 516672 3752 516724
rect 3700 516400 3752 516452
rect 9036 516400 9088 516452
rect 545028 516128 545080 516180
rect 546132 516128 546184 516180
rect 544660 511844 544712 511896
rect 545948 511844 546000 511896
rect 574100 509260 574152 509312
rect 577504 509260 577556 509312
rect 3608 507424 3660 507476
rect 3608 507220 3660 507272
rect 3516 507152 3568 507204
rect 7932 507152 7984 507204
rect 563796 507084 563848 507136
rect 574100 507084 574152 507136
rect 544660 506472 544712 506524
rect 554136 506472 554188 506524
rect 542084 505928 542136 505980
rect 542636 505928 542688 505980
rect 548708 503684 548760 503736
rect 579988 503684 580040 503736
rect 549352 501576 549404 501628
rect 580540 501576 580592 501628
rect 548800 500896 548852 500948
rect 579712 500896 579764 500948
rect 8852 499468 8904 499520
rect 38752 499468 38804 499520
rect 545028 498176 545080 498228
rect 547788 498176 547840 498228
rect 26884 494028 26936 494080
rect 38752 494028 38804 494080
rect 551652 494028 551704 494080
rect 579988 494028 580040 494080
rect 544660 493892 544712 493944
rect 549352 493892 549404 493944
rect 558920 492328 558972 492380
rect 563796 492328 563848 492380
rect 554044 489880 554096 489932
rect 580172 489880 580224 489932
rect 544660 489540 544712 489592
rect 545672 489540 545724 489592
rect 8024 488520 8076 488572
rect 38752 488520 38804 488572
rect 550824 488520 550876 488572
rect 558920 488520 558972 488572
rect 543372 485800 543424 485852
rect 545028 485800 545080 485852
rect 3516 485732 3568 485784
rect 38752 485732 38804 485784
rect 548800 484372 548852 484424
rect 580172 484372 580224 484424
rect 547512 478864 547564 478916
rect 579620 478864 579672 478916
rect 545948 474716 546000 474768
rect 580172 474716 580224 474768
rect 3516 471996 3568 472048
rect 10784 471996 10836 472048
rect 2964 471860 3016 471912
rect 3516 471860 3568 471912
rect 552940 469208 552992 469260
rect 579988 469208 580040 469260
rect 3148 467304 3200 467356
rect 7748 467304 7800 467356
rect 544660 466420 544712 466472
rect 561036 466420 561088 466472
rect 2964 463632 3016 463684
rect 38752 463632 38804 463684
rect 544660 462612 544712 462664
rect 548800 462612 548852 462664
rect 3148 462408 3200 462460
rect 7932 462408 7984 462460
rect 547604 460844 547656 460896
rect 580172 460844 580224 460896
rect 3056 459484 3108 459536
rect 38752 459484 38804 459536
rect 543464 458804 543516 458856
rect 562048 458804 562100 458856
rect 562048 455404 562100 455456
rect 566464 455404 566516 455456
rect 39948 455336 40000 455388
rect 41236 455336 41288 455388
rect 550088 454044 550140 454096
rect 580172 454044 580224 454096
rect 3240 452888 3292 452940
rect 9588 452888 9640 452940
rect 544660 452616 544712 452668
rect 574744 452616 574796 452668
rect 548800 449896 548852 449948
rect 580172 449896 580224 449948
rect 544660 449828 544712 449880
rect 580540 449828 580592 449880
rect 37464 449216 37516 449268
rect 39304 449216 39356 449268
rect 3148 447108 3200 447160
rect 13084 447108 13136 447160
rect 3240 444388 3292 444440
rect 38752 444388 38804 444440
rect 547604 444388 547656 444440
rect 580172 444388 580224 444440
rect 566464 442212 566516 442264
rect 574100 442212 574152 442264
rect 544936 440308 544988 440360
rect 550088 440308 550140 440360
rect 39488 440240 39540 440292
rect 41052 440240 41104 440292
rect 551744 440240 551796 440292
rect 580172 440240 580224 440292
rect 3240 438812 3292 438864
rect 11704 438812 11756 438864
rect 574100 437384 574152 437436
rect 577504 437384 577556 437436
rect 543924 435684 543976 435736
rect 545580 435684 545632 435736
rect 550088 434732 550140 434784
rect 580172 434732 580224 434784
rect 2964 431876 3016 431928
rect 38752 431876 38804 431928
rect 577504 431400 577556 431452
rect 579620 431400 579672 431452
rect 543924 431332 543976 431384
rect 545488 431332 545540 431384
rect 3240 429020 3292 429072
rect 6736 429020 6788 429072
rect 21456 426436 21508 426488
rect 38752 426436 38804 426488
rect 548892 425076 548944 425128
rect 580172 425076 580224 425128
rect 3240 423308 3292 423360
rect 9496 423308 9548 423360
rect 41052 418140 41104 418192
rect 41696 418140 41748 418192
rect 3240 418072 3292 418124
rect 9404 418072 9456 418124
rect 544200 417732 544252 417784
rect 546868 417732 546920 417784
rect 3148 413652 3200 413704
rect 6644 413652 6696 413704
rect 9588 412632 9640 412684
rect 38752 412632 38804 412684
rect 552572 409844 552624 409896
rect 580172 409844 580224 409896
rect 544200 409028 544252 409080
rect 546776 409028 546828 409080
rect 2780 408348 2832 408400
rect 5172 408348 5224 408400
rect 39396 405900 39448 405952
rect 41144 405900 41196 405952
rect 553124 405696 553176 405748
rect 580172 405696 580224 405748
rect 544936 405628 544988 405680
rect 552572 405628 552624 405680
rect 3240 404268 3292 404320
rect 29644 404268 29696 404320
rect 562324 401548 562376 401600
rect 579712 401548 579764 401600
rect 544844 400392 544896 400444
rect 544844 400188 544896 400240
rect 544752 400120 544804 400172
rect 553124 400120 553176 400172
rect 6828 398828 6880 398880
rect 38752 398828 38804 398880
rect 3240 398556 3292 398608
rect 9312 398556 9364 398608
rect 569868 398080 569920 398132
rect 580632 398080 580684 398132
rect 544936 397400 544988 397452
rect 550364 397400 550416 397452
rect 544752 395972 544804 396024
rect 551744 395972 551796 396024
rect 557540 395292 557592 395344
rect 569868 395292 569920 395344
rect 2780 393592 2832 393644
rect 5172 393592 5224 393644
rect 550364 391212 550416 391264
rect 563060 391212 563112 391264
rect 551192 390804 551244 390856
rect 557540 390804 557592 390856
rect 544752 390600 544804 390652
rect 551928 390600 551980 390652
rect 551744 390532 551796 390584
rect 579620 390532 579672 390584
rect 563060 388424 563112 388476
rect 570604 388424 570656 388476
rect 548984 386384 549036 386436
rect 580172 386384 580224 386436
rect 548340 386112 548392 386164
rect 551192 386112 551244 386164
rect 2780 384752 2832 384804
rect 5264 384752 5316 384804
rect 543188 382576 543240 382628
rect 550548 382576 550600 382628
rect 570604 382168 570656 382220
rect 579804 382168 579856 382220
rect 546040 380944 546092 380996
rect 548340 380944 548392 380996
rect 550548 378088 550600 378140
rect 552572 378088 552624 378140
rect 544752 377476 544804 377528
rect 550180 377476 550232 377528
rect 550272 376660 550324 376712
rect 580172 376660 580224 376712
rect 552572 374892 552624 374944
rect 558368 374892 558420 374944
rect 551836 372512 551888 372564
rect 579620 372512 579672 372564
rect 3240 368500 3292 368552
rect 33876 368500 33928 368552
rect 551836 365712 551888 365764
rect 580172 365712 580224 365764
rect 544752 364148 544804 364200
rect 545396 364148 545448 364200
rect 544844 362924 544896 362976
rect 545396 362924 545448 362976
rect 574836 361564 574888 361616
rect 580172 361564 580224 361616
rect 544936 358776 544988 358828
rect 560944 358776 560996 358828
rect 550180 356056 550232 356108
rect 579988 356056 580040 356108
rect 3148 354628 3200 354680
rect 10876 354628 10928 354680
rect 561036 353200 561088 353252
rect 580172 353200 580224 353252
rect 558276 352520 558328 352572
rect 574836 352520 574888 352572
rect 6644 350548 6696 350600
rect 38752 350548 38804 350600
rect 558368 350140 558420 350192
rect 561036 350140 561088 350192
rect 2780 349188 2832 349240
rect 5264 349188 5316 349240
rect 5356 346400 5408 346452
rect 38752 346400 38804 346452
rect 553308 346400 553360 346452
rect 580172 346400 580224 346452
rect 3332 344360 3384 344412
rect 9312 344360 9364 344412
rect 544752 342184 544804 342236
rect 553308 342184 553360 342236
rect 561036 340824 561088 340876
rect 569224 340824 569276 340876
rect 3332 339464 3384 339516
rect 9404 339464 9456 339516
rect 546132 338036 546184 338088
rect 580172 338036 580224 338088
rect 543004 336676 543056 336728
rect 546408 336676 546460 336728
rect 2964 334840 3016 334892
rect 6460 334840 6512 334892
rect 569224 334364 569276 334416
rect 574100 334364 574152 334416
rect 3332 332596 3384 332648
rect 38752 332596 38804 332648
rect 541900 330964 541952 331016
rect 547696 330964 547748 331016
rect 39580 329740 39632 329792
rect 40776 329740 40828 329792
rect 3240 328720 3292 328772
rect 6460 328720 6512 328772
rect 574100 328380 574152 328432
rect 579988 328380 580040 328432
rect 37096 324232 37148 324284
rect 38752 324232 38804 324284
rect 547696 322872 547748 322924
rect 579804 322872 579856 322924
rect 544936 318928 544988 318980
rect 550272 318928 550324 318980
rect 37464 318792 37516 318844
rect 39304 318792 39356 318844
rect 546132 316684 546184 316736
rect 558276 316684 558328 316736
rect 3332 315936 3384 315988
rect 26884 315936 26936 315988
rect 2964 314644 3016 314696
rect 38752 314644 38804 314696
rect 575480 313896 575532 313948
rect 580724 313896 580776 313948
rect 551928 313216 551980 313268
rect 580172 313216 580224 313268
rect 559656 311108 559708 311160
rect 575480 311108 575532 311160
rect 3332 310496 3384 310548
rect 38752 310496 38804 310548
rect 550272 307708 550324 307760
rect 580172 307708 580224 307760
rect 16488 306280 16540 306332
rect 38752 306280 38804 306332
rect 2780 304988 2832 305040
rect 5356 304988 5408 305040
rect 556160 302336 556212 302388
rect 559656 302336 559708 302388
rect 577504 302268 577556 302320
rect 580816 302268 580868 302320
rect 550272 302200 550324 302252
rect 580172 302200 580224 302252
rect 553124 299548 553176 299600
rect 556160 299548 556212 299600
rect 550364 296692 550416 296744
rect 579620 296692 579672 296744
rect 3332 295264 3384 295316
rect 21456 295264 21508 295316
rect 35164 293904 35216 293956
rect 38752 293904 38804 293956
rect 547696 292544 547748 292596
rect 579804 292544 579856 292596
rect 3148 289824 3200 289876
rect 11704 289824 11756 289876
rect 546224 287648 546276 287700
rect 553124 287648 553176 287700
rect 563336 287648 563388 287700
rect 577504 287648 577556 287700
rect 550548 287036 550600 287088
rect 579620 287036 579672 287088
rect 561036 284316 561088 284368
rect 563336 284316 563388 284368
rect 14464 284248 14516 284300
rect 38752 284248 38804 284300
rect 547788 284248 547840 284300
rect 579620 284248 579672 284300
rect 3332 280440 3384 280492
rect 9496 280440 9548 280492
rect 37556 280100 37608 280152
rect 39304 280100 39356 280152
rect 544936 278740 544988 278792
rect 553308 278740 553360 278792
rect 553032 278672 553084 278724
rect 579988 278672 580040 278724
rect 544752 275612 544804 275664
rect 550456 275612 550508 275664
rect 39396 275340 39448 275392
rect 40868 275340 40920 275392
rect 3332 274660 3384 274712
rect 10876 274660 10928 274712
rect 553308 274592 553360 274644
rect 580172 274592 580224 274644
rect 554780 273912 554832 273964
rect 561036 273912 561088 273964
rect 553032 270716 553084 270768
rect 554780 270716 554832 270768
rect 6552 270444 6604 270496
rect 38752 270444 38804 270496
rect 546316 266976 546368 267028
rect 553032 266976 553084 267028
rect 3148 266092 3200 266144
rect 9588 266092 9640 266144
rect 546408 265684 546460 265736
rect 556896 265684 556948 265736
rect 547052 265616 547104 265668
rect 563060 265616 563112 265668
rect 3148 260176 3200 260228
rect 9588 260176 9640 260228
rect 563060 260108 563112 260160
rect 579804 260108 579856 260160
rect 551928 258068 551980 258120
rect 580172 258068 580224 258120
rect 544752 255280 544804 255332
rect 550456 255280 550508 255332
rect 556896 251812 556948 251864
rect 572720 251812 572772 251864
rect 37556 251200 37608 251252
rect 38752 251200 38804 251252
rect 572720 249704 572772 249756
rect 579620 249704 579672 249756
rect 37648 248072 37700 248124
rect 38844 248072 38896 248124
rect 544752 247052 544804 247104
rect 553032 247052 553084 247104
rect 3608 246100 3660 246152
rect 8116 246100 8168 246152
rect 11704 244196 11756 244248
rect 38752 244196 38804 244248
rect 544752 242904 544804 242956
rect 561036 242904 561088 242956
rect 3608 241068 3660 241120
rect 9128 241068 9180 241120
rect 37740 240048 37792 240100
rect 38752 240048 38804 240100
rect 545672 240048 545724 240100
rect 580172 240048 580224 240100
rect 544752 237396 544804 237448
rect 551192 237396 551244 237448
rect 3608 236172 3660 236224
rect 7840 236172 7892 236224
rect 21364 234540 21416 234592
rect 38752 234540 38804 234592
rect 553032 234540 553084 234592
rect 579988 234540 580040 234592
rect 544476 229780 544528 229832
rect 547420 229780 547472 229832
rect 574008 229100 574060 229152
rect 580172 229100 580224 229152
rect 3148 226312 3200 226364
rect 6552 226312 6604 226364
rect 544752 224952 544804 225004
rect 553124 224952 553176 225004
rect 570604 223252 570656 223304
rect 574008 223252 574060 223304
rect 3148 220804 3200 220856
rect 38844 220804 38896 220856
rect 544752 219444 544804 219496
rect 553032 219444 553084 219496
rect 560944 219376 560996 219428
rect 579804 219376 579856 219428
rect 574744 215228 574796 215280
rect 580172 215228 580224 215280
rect 3608 212440 3660 212492
rect 33784 212440 33836 212492
rect 3056 211284 3108 211336
rect 3608 211284 3660 211336
rect 544476 211148 544528 211200
rect 547420 211148 547472 211200
rect 553124 209720 553176 209772
rect 579988 209720 580040 209772
rect 553400 209040 553452 209092
rect 570604 209040 570656 209092
rect 9220 208292 9272 208344
rect 38844 208292 38896 208344
rect 544752 208292 544804 208344
rect 564440 208292 564492 208344
rect 551100 205640 551152 205692
rect 553400 205640 553452 205692
rect 3884 201424 3936 201476
rect 5448 201424 5500 201476
rect 553032 200064 553084 200116
rect 580172 200064 580224 200116
rect 3148 196664 3200 196716
rect 9128 196664 9180 196716
rect 549076 195984 549128 196036
rect 551100 195984 551152 196036
rect 5448 194488 5500 194540
rect 8116 194488 8168 194540
rect 547420 194488 547472 194540
rect 580172 194488 580224 194540
rect 11704 193196 11756 193248
rect 38844 193196 38896 193248
rect 554136 190408 554188 190460
rect 579620 190408 579672 190460
rect 37832 190068 37884 190120
rect 39488 190068 39540 190120
rect 544476 189524 544528 189576
rect 546408 189524 546460 189576
rect 3148 186600 3200 186652
rect 7840 186600 7892 186652
rect 3056 184900 3108 184952
rect 38844 184900 38896 184952
rect 546408 184900 546460 184952
rect 549812 184832 549864 184884
rect 552848 184832 552900 184884
rect 580172 184832 580224 184884
rect 544752 183540 544804 183592
rect 565084 183540 565136 183592
rect 3148 182112 3200 182164
rect 10692 182112 10744 182164
rect 546408 180820 546460 180872
rect 549076 180820 549128 180872
rect 548616 180752 548668 180804
rect 579988 180752 580040 180804
rect 543832 180548 543884 180600
rect 546684 180548 546736 180600
rect 549812 178032 549864 178084
rect 554688 177964 554740 178016
rect 3056 176944 3108 176996
rect 6736 176944 6788 176996
rect 13084 176604 13136 176656
rect 38844 176604 38896 176656
rect 544752 176604 544804 176656
rect 559564 176604 559616 176656
rect 550456 175176 550508 175228
rect 579620 175176 579672 175228
rect 8116 173816 8168 173868
rect 12072 173816 12124 173868
rect 554780 172932 554832 172984
rect 558920 172932 558972 172984
rect 3884 172456 3936 172508
rect 5448 172456 5500 172508
rect 3056 172116 3108 172168
rect 9220 172116 9272 172168
rect 545672 171776 545724 171828
rect 580908 171776 580960 171828
rect 544476 171232 544528 171284
rect 547420 171232 547472 171284
rect 558920 170348 558972 170400
rect 569684 170348 569736 170400
rect 9588 168308 9640 168360
rect 38844 168308 38896 168360
rect 543832 167220 543884 167272
rect 546592 167220 546644 167272
rect 569684 167016 569736 167068
rect 574744 166948 574796 167000
rect 12072 166540 12124 166592
rect 14464 166540 14516 166592
rect 5448 165520 5500 165572
rect 8116 165520 8168 165572
rect 547788 164228 547840 164280
rect 579988 164228 580040 164280
rect 2780 162460 2832 162512
rect 5080 162460 5132 162512
rect 17868 161440 17920 161492
rect 38844 161440 38896 161492
rect 574744 160080 574796 160132
rect 580172 160012 580224 160064
rect 544752 158652 544804 158704
rect 556804 158652 556856 158704
rect 14464 155864 14516 155916
rect 15200 155864 15252 155916
rect 565084 155864 565136 155916
rect 579620 155864 579672 155916
rect 3792 153144 3844 153196
rect 5356 153144 5408 153196
rect 15200 152056 15252 152108
rect 17224 152056 17276 152108
rect 548616 149064 548668 149116
rect 579620 149064 579672 149116
rect 3424 147568 3476 147620
rect 25504 147568 25556 147620
rect 8116 144848 8168 144900
rect 11796 144848 11848 144900
rect 17224 144848 17276 144900
rect 18052 144848 18104 144900
rect 2780 142332 2832 142384
rect 5080 142332 5132 142384
rect 18052 141108 18104 141160
rect 21180 141108 21232 141160
rect 547328 140700 547380 140752
rect 580172 140700 580224 140752
rect 5540 140292 5592 140344
rect 8208 140292 8260 140344
rect 39948 139476 40000 139528
rect 40960 139476 41012 139528
rect 3608 139408 3660 139460
rect 21180 139408 21232 139460
rect 6092 139340 6144 139392
rect 24216 139340 24268 139392
rect 8208 137844 8260 137896
rect 9588 137844 9640 137896
rect 3424 137504 3476 137556
rect 8116 137504 8168 137556
rect 11796 137504 11848 137556
rect 14464 137504 14516 137556
rect 549076 135260 549128 135312
rect 579620 135260 579672 135312
rect 33876 132404 33928 132456
rect 38844 132404 38896 132456
rect 24216 131112 24268 131164
rect 25504 131112 25556 131164
rect 6092 131044 6144 131096
rect 8852 131044 8904 131096
rect 551192 131044 551244 131096
rect 579804 131044 579856 131096
rect 3240 128256 3292 128308
rect 10600 128256 10652 128308
rect 8852 126896 8904 126948
rect 13084 126896 13136 126948
rect 14464 126896 14516 126948
rect 15200 126896 15252 126948
rect 9588 126828 9640 126880
rect 15844 126828 15896 126880
rect 3148 125604 3200 125656
rect 3700 125536 3752 125588
rect 4712 125536 4764 125588
rect 5540 125536 5592 125588
rect 15200 123156 15252 123208
rect 17224 123156 17276 123208
rect 3608 122952 3660 123004
rect 8208 122952 8260 123004
rect 13084 122204 13136 122256
rect 14372 122204 14424 122256
rect 5540 120980 5592 121032
rect 7472 120980 7524 121032
rect 552848 120096 552900 120148
rect 580172 120096 580224 120148
rect 4712 118600 4764 118652
rect 5540 118600 5592 118652
rect 3608 117308 3660 117360
rect 12440 117308 12492 117360
rect 14372 117240 14424 117292
rect 17316 117240 17368 117292
rect 561036 117240 561088 117292
rect 579620 117240 579672 117292
rect 7472 117036 7524 117088
rect 9588 117036 9640 117088
rect 12440 115744 12492 115796
rect 16212 115744 16264 115796
rect 5540 115608 5592 115660
rect 7472 115608 7524 115660
rect 25504 115132 25556 115184
rect 27620 115132 27672 115184
rect 20628 114452 20680 114504
rect 38844 114452 38896 114504
rect 544660 114452 544712 114504
rect 558184 114452 558236 114504
rect 3056 113160 3108 113212
rect 6092 113160 6144 113212
rect 9588 110440 9640 110492
rect 17316 110440 17368 110492
rect 12440 110372 12492 110424
rect 27620 110440 27672 110492
rect 29644 110440 29696 110492
rect 567752 110440 567804 110492
rect 580172 110440 580224 110492
rect 20168 110372 20220 110424
rect 7472 109624 7524 109676
rect 10600 109624 10652 109676
rect 3332 109556 3384 109608
rect 5356 109556 5408 109608
rect 10784 108944 10836 108996
rect 38844 108944 38896 108996
rect 3148 108672 3200 108724
rect 6644 108672 6696 108724
rect 16212 108264 16264 108316
rect 19984 108264 20036 108316
rect 5356 107584 5408 107636
rect 6644 107584 6696 107636
rect 12440 107584 12492 107636
rect 17408 107584 17460 107636
rect 20168 107584 20220 107636
rect 22836 107584 22888 107636
rect 17224 107516 17276 107568
rect 20076 107516 20128 107568
rect 17408 104796 17460 104848
rect 18328 104796 18380 104848
rect 543556 104116 543608 104168
rect 567752 104116 567804 104168
rect 3332 103436 3384 103488
rect 24124 103436 24176 103488
rect 6644 102620 6696 102672
rect 7472 102620 7524 102672
rect 20076 102484 20128 102536
rect 21548 102484 21600 102536
rect 578240 102144 578292 102196
rect 580172 102144 580224 102196
rect 549996 102076 550048 102128
rect 579620 102076 579672 102128
rect 18328 100988 18380 101040
rect 21364 100988 21416 101040
rect 19984 100716 20036 100768
rect 21456 100716 21508 100768
rect 21548 100580 21600 100632
rect 22744 100580 22796 100632
rect 15844 99968 15896 100020
rect 20720 99968 20772 100020
rect 22836 99084 22888 99136
rect 24124 99084 24176 99136
rect 7472 99016 7524 99068
rect 8852 99016 8904 99068
rect 10600 98812 10652 98864
rect 11796 98812 11848 98864
rect 39120 97928 39172 97980
rect 41144 97928 41196 97980
rect 566464 97248 566516 97300
rect 578148 97248 578200 97300
rect 8852 96568 8904 96620
rect 16488 96568 16540 96620
rect 20720 95140 20772 95192
rect 22836 95140 22888 95192
rect 543372 95140 543424 95192
rect 543740 95140 543792 95192
rect 563796 94460 563848 94512
rect 580724 94460 580776 94512
rect 40960 93508 41012 93560
rect 41604 93508 41656 93560
rect 2780 92760 2832 92812
rect 5356 92760 5408 92812
rect 16580 92488 16632 92540
rect 25688 92420 25740 92472
rect 38936 92012 38988 92064
rect 41052 92012 41104 92064
rect 11796 91876 11848 91928
rect 13728 91876 13780 91928
rect 22744 91060 22796 91112
rect 25504 90992 25556 91044
rect 561772 89700 561824 89752
rect 566464 89700 566516 89752
rect 13728 88340 13780 88392
rect 15200 88272 15252 88324
rect 24124 88272 24176 88324
rect 25596 88272 25648 88324
rect 29644 88272 29696 88324
rect 32404 88272 32456 88324
rect 22836 86912 22888 86964
rect 24124 86912 24176 86964
rect 544844 86232 544896 86284
rect 563796 86232 563848 86284
rect 15200 85552 15252 85604
rect 558828 85552 558880 85604
rect 561772 85552 561824 85604
rect 18604 85484 18656 85536
rect 21456 84192 21508 84244
rect 551192 84192 551244 84244
rect 558828 84192 558880 84244
rect 23940 84124 23992 84176
rect 25688 83104 25740 83156
rect 27528 83104 27580 83156
rect 3332 82832 3384 82884
rect 24860 82764 24912 82816
rect 39856 82628 39908 82680
rect 41328 82628 41380 82680
rect 40040 82356 40092 82408
rect 41512 82356 41564 82408
rect 543832 81404 543884 81456
rect 558184 81404 558236 81456
rect 545764 81336 545816 81388
rect 580172 81336 580224 81388
rect 549536 79772 549588 79824
rect 551192 79772 551244 79824
rect 23940 79364 23992 79416
rect 25780 79364 25832 79416
rect 27528 79024 27580 79076
rect 29000 79024 29052 79076
rect 2780 78684 2832 78736
rect 5448 78684 5500 78736
rect 24860 78616 24912 78668
rect 27252 78616 27304 78668
rect 32404 78616 32456 78668
rect 36544 78616 36596 78668
rect 21364 77256 21416 77308
rect 18604 77188 18656 77240
rect 20628 77188 20680 77240
rect 29000 77256 29052 77308
rect 25412 77188 25464 77240
rect 33784 77188 33836 77240
rect 25504 77052 25556 77104
rect 26976 77052 27028 77104
rect 25596 75896 25648 75948
rect 26884 75896 26936 75948
rect 27252 75828 27304 75880
rect 30288 75828 30340 75880
rect 543648 75828 543700 75880
rect 549536 75896 549588 75948
rect 24124 74536 24176 74588
rect 3332 74468 3384 74520
rect 10416 74468 10468 74520
rect 27528 74468 27580 74520
rect 39948 73652 40000 73704
rect 41696 73652 41748 73704
rect 542268 73176 542320 73228
rect 543556 73176 543608 73228
rect 25780 73108 25832 73160
rect 27252 73108 27304 73160
rect 27528 71748 27580 71800
rect 29092 71680 29144 71732
rect 27252 70456 27304 70508
rect 31024 70456 31076 70508
rect 30380 69844 30432 69896
rect 35164 69844 35216 69896
rect 25412 69028 25464 69080
rect 29092 69028 29144 69080
rect 27620 68960 27672 69012
rect 32496 68960 32548 69012
rect 543832 68960 543884 69012
rect 554044 68960 554096 69012
rect 3332 68892 3384 68944
rect 8024 68892 8076 68944
rect 20720 68280 20772 68332
rect 29644 68280 29696 68332
rect 27620 67532 27672 67584
rect 30288 67532 30340 67584
rect 575480 66240 575532 66292
rect 578976 66240 579028 66292
rect 38844 64744 38896 64796
rect 40960 64744 41012 64796
rect 31024 64132 31076 64184
rect 32404 64132 32456 64184
rect 543832 64132 543884 64184
rect 545948 64132 546000 64184
rect 2780 63996 2832 64048
rect 4804 63996 4856 64048
rect 26976 63724 27028 63776
rect 31484 63724 31536 63776
rect 35164 63520 35216 63572
rect 38108 63452 38160 63504
rect 30288 62636 30340 62688
rect 32312 62636 32364 62688
rect 571708 62024 571760 62076
rect 575388 62092 575440 62144
rect 33784 60596 33836 60648
rect 34520 60596 34572 60648
rect 26884 60188 26936 60240
rect 31668 60188 31720 60240
rect 543832 59508 543884 59560
rect 546500 59508 546552 59560
rect 3700 59372 3752 59424
rect 38844 59372 38896 59424
rect 31484 59304 31536 59356
rect 33140 59304 33192 59356
rect 567936 59304 567988 59356
rect 571708 59304 571760 59356
rect 32312 57876 32364 57928
rect 34428 57876 34480 57928
rect 31760 56584 31812 56636
rect 35624 56516 35676 56568
rect 39212 56516 39264 56568
rect 41236 56516 41288 56568
rect 33140 56108 33192 56160
rect 36636 56108 36688 56160
rect 34520 55700 34572 55752
rect 36820 55700 36872 55752
rect 543832 53796 543884 53848
rect 35624 53048 35676 53100
rect 41420 53048 41472 53100
rect 564440 52776 564492 52828
rect 567936 52776 567988 52828
rect 38108 52436 38160 52488
rect 39212 52436 39264 52488
rect 567844 52368 567896 52420
rect 579988 52368 580040 52420
rect 32496 52300 32548 52352
rect 36728 52300 36780 52352
rect 29644 51620 29696 51672
rect 34428 51620 34480 51672
rect 36820 51348 36872 51400
rect 38108 51348 38160 51400
rect 41420 50847 41472 50856
rect 41420 50813 41429 50847
rect 41429 50813 41463 50847
rect 41463 50813 41472 50847
rect 41420 50804 41472 50813
rect 40960 50668 41012 50720
rect 41420 50668 41472 50720
rect 40316 50600 40368 50652
rect 40316 50464 40368 50516
rect 40592 50464 40644 50516
rect 40500 50260 40552 50312
rect 34520 49716 34572 49768
rect 38200 49648 38252 49700
rect 2780 48288 2832 48340
rect 4712 48288 4764 48340
rect 34520 47608 34572 47660
rect 36268 47608 36320 47660
rect 559840 47472 559892 47524
rect 564440 47472 564492 47524
rect 544660 46971 544712 46980
rect 544660 46937 544669 46971
rect 544669 46937 544703 46971
rect 544703 46937 544712 46971
rect 544660 46928 544712 46937
rect 32404 46860 32456 46912
rect 34520 46860 34572 46912
rect 36636 46860 36688 46912
rect 37280 46860 37332 46912
rect 551560 46860 551612 46912
rect 579988 46860 580040 46912
rect 544660 46792 544712 46844
rect 563704 46792 563756 46844
rect 544660 46044 544712 46096
rect 544844 46044 544896 46096
rect 544844 45908 544896 45960
rect 545028 45908 545080 45960
rect 41788 45815 41840 45824
rect 41788 45781 41797 45815
rect 41797 45781 41831 45815
rect 41831 45781 41840 45815
rect 41788 45772 41840 45781
rect 545028 45772 545080 45824
rect 41420 45704 41472 45756
rect 40500 45568 40552 45620
rect 41420 45611 41472 45620
rect 41420 45577 41429 45611
rect 41429 45577 41463 45611
rect 41463 45577 41472 45611
rect 41420 45568 41472 45577
rect 41880 45514 41932 45566
rect 552020 45500 552072 45552
rect 559840 45568 559892 45620
rect 36268 44956 36320 45008
rect 38844 44956 38896 45008
rect 3240 44752 3292 44804
rect 3516 44752 3568 44804
rect 580540 44752 580592 44804
rect 580724 44752 580776 44804
rect 37096 44616 37148 44668
rect 542820 44659 542872 44668
rect 542820 44625 542829 44659
rect 542829 44625 542863 44659
rect 542863 44625 542872 44659
rect 542820 44616 542872 44625
rect 37556 44548 37608 44600
rect 580908 44548 580960 44600
rect 3608 44480 3660 44532
rect 3792 44480 3844 44532
rect 40592 44480 40644 44532
rect 580080 44480 580132 44532
rect 38200 44412 38252 44464
rect 40592 44387 40644 44396
rect 40592 44353 40601 44387
rect 40601 44353 40635 44387
rect 40635 44353 40644 44387
rect 40592 44344 40644 44353
rect 40960 44412 41012 44464
rect 580448 44412 580500 44464
rect 544936 44344 544988 44396
rect 34428 44276 34480 44328
rect 543648 44276 543700 44328
rect 39212 44208 39264 44260
rect 542176 44208 542228 44260
rect 542820 44208 542872 44260
rect 544476 44208 544528 44260
rect 39028 44140 39080 44192
rect 40960 44140 41012 44192
rect 41880 44183 41932 44192
rect 41880 44149 41889 44183
rect 41889 44149 41923 44183
rect 41923 44149 41932 44183
rect 41880 44140 41932 44149
rect 543372 44140 543424 44192
rect 543556 44140 543608 44192
rect 544752 44140 544804 44192
rect 34520 44072 34572 44124
rect 544200 44072 544252 44124
rect 36544 44004 36596 44056
rect 543924 44004 543976 44056
rect 39304 43936 39356 43988
rect 39672 43868 39724 43920
rect 542176 43936 542228 43988
rect 38752 43800 38804 43852
rect 546132 43868 546184 43920
rect 546408 43800 546460 43852
rect 39764 43732 39816 43784
rect 546040 43732 546092 43784
rect 36728 43664 36780 43716
rect 542728 43664 542780 43716
rect 41604 43596 41656 43648
rect 546316 43596 546368 43648
rect 37280 43528 37332 43580
rect 541900 43528 541952 43580
rect 542728 43528 542780 43580
rect 20628 43460 20680 43512
rect 544844 43460 544896 43512
rect 4804 43392 4856 43444
rect 544292 43392 544344 43444
rect 41512 43324 41564 43376
rect 544660 43324 544712 43376
rect 41880 43256 41932 43308
rect 542820 43256 542872 43308
rect 41144 43188 41196 43240
rect 542268 43188 542320 43240
rect 41328 43120 41380 43172
rect 546224 43120 546276 43172
rect 41420 43052 41472 43104
rect 542176 43052 542228 43104
rect 41880 42984 41932 43036
rect 558184 42712 558236 42764
rect 580172 42712 580224 42764
rect 545304 42576 545356 42628
rect 543280 42508 543332 42560
rect 40316 42440 40368 42492
rect 543740 42440 543792 42492
rect 40132 42372 40184 42424
rect 196072 42372 196124 42424
rect 379428 42372 379480 42424
rect 542452 42372 542504 42424
rect 38936 42304 38988 42356
rect 231860 42304 231912 42356
rect 277308 42304 277360 42356
rect 545028 42304 545080 42356
rect 4160 42236 4212 42288
rect 320180 42236 320232 42288
rect 333888 42236 333940 42288
rect 543832 42236 543884 42288
rect 40592 42168 40644 42220
rect 382280 42168 382332 42220
rect 395988 42168 396040 42220
rect 543464 42168 543516 42220
rect 169668 42100 169720 42152
rect 544384 42100 544436 42152
rect 39948 42032 40000 42084
rect 580448 42032 580500 42084
rect 191840 42007 191892 42016
rect 191840 41973 191849 42007
rect 191849 41973 191883 42007
rect 191883 41973 191892 42007
rect 191840 41964 191892 41973
rect 436008 42007 436060 42016
rect 436008 41973 436017 42007
rect 436017 41973 436051 42007
rect 436051 41973 436060 42007
rect 436008 41964 436060 41973
rect 509148 42007 509200 42016
rect 509148 41973 509157 42007
rect 509157 41973 509191 42007
rect 509191 41973 509200 42007
rect 509148 41964 509200 41973
rect 536748 42007 536800 42016
rect 536748 41973 536757 42007
rect 536757 41973 536791 42007
rect 536791 41973 536800 42007
rect 536748 41964 536800 41973
rect 538312 41420 538364 41472
rect 542360 41420 542412 41472
rect 3332 41352 3384 41404
rect 65984 41352 66036 41404
rect 157432 41352 157484 41404
rect 162860 41352 162912 41404
rect 384672 41352 384724 41404
rect 547696 41352 547748 41404
rect 7840 41284 7892 41336
rect 71780 41284 71832 41336
rect 305920 41284 305972 41336
rect 547788 41284 547840 41336
rect 7564 41216 7616 41268
rect 156604 41216 156656 41268
rect 275560 41216 275612 41268
rect 547236 41216 547288 41268
rect 33048 41148 33100 41200
rect 329196 41148 329248 41200
rect 366456 41148 366508 41200
rect 552756 41148 552808 41200
rect 9128 41080 9180 41132
rect 168748 41080 168800 41132
rect 245200 41080 245252 41132
rect 548524 41080 548576 41132
rect 5264 41012 5316 41064
rect 226340 41012 226392 41064
rect 269488 41012 269540 41064
rect 580356 41012 580408 41064
rect 4896 40944 4948 40996
rect 232780 40944 232832 40996
rect 238760 40944 238812 40996
rect 571340 40944 571392 40996
rect 7748 40876 7800 40928
rect 347780 40876 347832 40928
rect 351000 40876 351052 40928
rect 548984 40876 549036 40928
rect 6552 40808 6604 40860
rect 408316 40808 408368 40860
rect 3424 40740 3476 40792
rect 411444 40740 411496 40792
rect 5356 40672 5408 40724
rect 420460 40672 420512 40724
rect 513288 40672 513340 40724
rect 542728 40672 542780 40724
rect 4712 40604 4764 40656
rect 69204 40604 69256 40656
rect 150992 40604 151044 40656
rect 580816 40604 580868 40656
rect 9036 40536 9088 40588
rect 441620 40536 441672 40588
rect 493232 40536 493284 40588
rect 545856 40536 545908 40588
rect 68008 40468 68060 40520
rect 135812 40468 135864 40520
rect 138848 40468 138900 40520
rect 580632 40468 580684 40520
rect 7932 40400 7984 40452
rect 96436 40400 96488 40452
rect 102600 40400 102652 40452
rect 547512 40400 547564 40452
rect 3976 40332 4028 40384
rect 465908 40332 465960 40384
rect 469128 40332 469180 40384
rect 580080 40332 580132 40384
rect 5080 40264 5132 40316
rect 474924 40264 474976 40316
rect 496360 40264 496412 40316
rect 580540 40264 580592 40316
rect 5448 40196 5500 40248
rect 499212 40196 499264 40248
rect 3792 40128 3844 40180
rect 508412 40128 508464 40180
rect 6736 40060 6788 40112
rect 520372 40060 520424 40112
rect 37188 39992 37240 40044
rect 51080 39992 51132 40044
rect 123760 39992 123812 40044
rect 345664 39992 345716 40044
rect 348240 39992 348292 40044
rect 352380 39992 352432 40044
rect 354956 39992 355008 40044
rect 511448 39992 511500 40044
rect 548892 39992 548944 40044
rect 41788 39924 41840 39976
rect 159916 39924 159968 39976
rect 314568 39924 314620 39976
rect 316040 39924 316092 39976
rect 529664 39924 529716 39976
rect 552940 39924 552992 39976
rect 5172 39856 5224 39908
rect 429660 39856 429712 39908
rect 535736 39856 535788 39908
rect 551468 39856 551520 39908
rect 3608 39788 3660 39840
rect 417516 39788 417568 39840
rect 426624 39788 426676 39840
rect 439504 39788 439556 39840
rect 450912 39788 450964 39840
rect 548800 39788 548852 39840
rect 1308 39720 1360 39772
rect 41972 39720 42024 39772
rect 65984 39720 66036 39772
rect 453764 39720 453816 39772
rect 459928 39720 459980 39772
rect 547604 39720 547656 39772
rect 2780 39652 2832 39704
rect 4988 39652 5040 39704
rect 9496 39652 9548 39704
rect 196348 39652 196400 39704
rect 208584 39652 208636 39704
rect 551928 39652 551980 39704
rect 9220 39584 9272 39636
rect 190276 39584 190328 39636
rect 211528 39584 211580 39636
rect 549076 39584 549128 39636
rect 8208 39516 8260 39568
rect 214564 39516 214616 39568
rect 217600 39516 217652 39568
rect 550364 39516 550416 39568
rect 9312 39448 9364 39500
rect 338764 39448 338816 39500
rect 344928 39448 344980 39500
rect 550088 39448 550140 39500
rect 8116 39380 8168 39432
rect 335636 39380 335688 39432
rect 369032 39380 369084 39432
rect 551744 39380 551796 39432
rect 13728 39312 13780 39364
rect 53932 39312 53984 39364
rect 59360 39312 59412 39364
rect 61384 39312 61436 39364
rect 86868 39312 86920 39364
rect 117596 39312 117648 39364
rect 126704 39312 126756 39364
rect 443644 39312 443696 39364
rect 514392 39312 514444 39364
rect 580264 39312 580316 39364
rect 6092 39244 6144 39296
rect 302332 39244 302384 39296
rect 332784 39244 332836 39296
rect 367744 39244 367796 39296
rect 375104 39244 375156 39296
rect 385040 39244 385092 39296
rect 387248 39244 387300 39296
rect 549904 39244 549956 39296
rect 9404 39176 9456 39228
rect 250812 39176 250864 39228
rect 260104 39176 260156 39228
rect 10876 39108 10928 39160
rect 241796 39108 241848 39160
rect 247960 39108 248012 39160
rect 259460 39108 259512 39160
rect 281264 39108 281316 39160
rect 551836 39108 551888 39160
rect 3516 39040 3568 39092
rect 178132 39040 178184 39092
rect 205456 39040 205508 39092
rect 285680 39040 285732 39092
rect 290280 39040 290332 39092
rect 548616 39040 548668 39092
rect 38384 38972 38436 39024
rect 181260 38972 181312 39024
rect 272248 38972 272300 39024
rect 301504 38972 301556 39024
rect 362960 38972 363012 39024
rect 372620 38972 372672 39024
rect 435640 38972 435692 39024
rect 451924 38972 451976 39024
rect 490288 38972 490340 39024
rect 548708 38972 548760 39024
rect 44088 38904 44140 38956
rect 81164 38904 81216 38956
rect 105544 38904 105596 38956
rect 159364 38904 159416 38956
rect 266268 38904 266320 38956
rect 293316 38904 293368 38956
rect 502432 38904 502484 38956
rect 547880 38904 547932 38956
rect 38292 38836 38344 38888
rect 47860 38836 47912 38888
rect 90456 38836 90508 38888
rect 131764 38836 131816 38888
rect 131856 38836 131908 38888
rect 172060 38836 172112 38888
rect 444840 38836 444892 38888
rect 6460 38768 6512 38820
rect 114652 38768 114704 38820
rect 119988 38768 120040 38820
rect 144920 38768 144972 38820
rect 154120 38768 154172 38820
rect 182824 38768 182876 38820
rect 254032 38768 254084 38820
rect 255228 38768 255280 38820
rect 414480 38768 414532 38820
rect 415308 38768 415360 38820
rect 482928 38768 482980 38820
rect 484124 38768 484176 38820
rect 538680 38768 538732 38820
rect 539508 38768 539560 38820
rect 541808 38836 541860 38888
rect 542268 38836 542320 38888
rect 550548 38836 550600 38888
rect 550180 38768 550232 38820
rect 41880 38700 41932 38752
rect 75276 38700 75328 38752
rect 129832 38700 129884 38752
rect 131028 38700 131080 38752
rect 550272 38700 550324 38752
rect 7656 38632 7708 38684
rect 44916 38632 44968 38684
rect 108672 38632 108724 38684
rect 552848 38632 552900 38684
rect 346308 38292 346360 38344
rect 350540 38292 350592 38344
rect 349988 37884 350040 37936
rect 352380 37884 352432 37936
rect 449808 37884 449860 37936
rect 544568 37884 544620 37936
rect 547144 37204 547196 37256
rect 580172 37204 580224 37256
rect 39488 36524 39540 36576
rect 368480 36524 368532 36576
rect 343548 35912 343600 35964
rect 346308 35912 346360 35964
rect 343640 35232 343692 35284
rect 349988 35232 350040 35284
rect 40040 35164 40092 35216
rect 349160 35164 349212 35216
rect 340512 34416 340564 34468
rect 345664 34484 345716 34536
rect 3424 34348 3476 34400
rect 8944 34348 8996 34400
rect 341524 33124 341576 33176
rect 343548 33124 343600 33176
rect 438768 33056 438820 33108
rect 580080 33056 580132 33108
rect 336004 31696 336056 31748
rect 340512 31764 340564 31816
rect 339684 31696 339736 31748
rect 343640 31764 343692 31816
rect 279424 31016 279476 31068
rect 287704 31016 287756 31068
rect 338028 29792 338080 29844
rect 339684 29792 339736 29844
rect 332600 27616 332652 27668
rect 338028 27616 338080 27668
rect 551376 27548 551428 27600
rect 580080 27548 580132 27600
rect 39580 25508 39632 25560
rect 498200 25508 498252 25560
rect 331220 25304 331272 25356
rect 336004 25304 336056 25356
rect 3240 24692 3292 24744
rect 6368 24692 6420 24744
rect 326620 23536 326672 23588
rect 331220 23536 331272 23588
rect 329840 23468 329892 23520
rect 332600 23468 332652 23520
rect 320824 22040 320876 22092
rect 326620 22108 326672 22160
rect 269120 19932 269172 19984
rect 279424 19932 279476 19984
rect 61384 17892 61436 17944
rect 64512 17892 64564 17944
rect 3424 15104 3476 15156
rect 11704 15104 11756 15156
rect 326344 15104 326396 15156
rect 329472 15172 329524 15224
rect 340144 15172 340196 15224
rect 341524 15172 341576 15224
rect 64512 10276 64564 10328
rect 69664 10276 69716 10328
rect 2964 9868 3016 9920
rect 6276 9868 6328 9920
rect 266176 8236 266228 8288
rect 580172 8236 580224 8288
rect 376116 6264 376168 6316
rect 545120 6264 545172 6316
rect 136364 6196 136416 6248
rect 456800 6196 456852 6248
rect 93124 6128 93176 6180
rect 542084 6128 542136 6180
rect 57888 5448 57940 5500
rect 242900 5448 242952 5500
rect 282828 5448 282880 5500
rect 544016 5448 544068 5500
rect 39856 5380 39908 5432
rect 352748 5380 352800 5432
rect 356060 5380 356112 5432
rect 545672 5380 545724 5432
rect 69756 5312 69808 5364
rect 186320 5312 186372 5364
rect 229652 5312 229704 5364
rect 542912 5312 542964 5364
rect 2780 5244 2832 5296
rect 4804 5244 4856 5296
rect 79876 5244 79928 5296
rect 396080 5244 396132 5296
rect 406108 5244 406160 5296
rect 545488 5244 545540 5296
rect 37924 5176 37976 5228
rect 409420 5176 409472 5228
rect 142988 5108 143040 5160
rect 544108 5108 544160 5160
rect 39396 5040 39448 5092
rect 452660 5040 452712 5092
rect 69664 4972 69716 5024
rect 126428 4972 126480 5024
rect 129740 4972 129792 5024
rect 545580 4972 545632 5024
rect 26516 4904 26568 4956
rect 480260 4904 480312 4956
rect 49884 4836 49936 4888
rect 541992 4836 542044 4888
rect 37464 4768 37516 4820
rect 542452 4768 542504 4820
rect 111708 4700 111760 4752
rect 256332 4700 256384 4752
rect 296260 4700 296312 4752
rect 340144 4700 340196 4752
rect 389364 4700 389416 4752
rect 505100 4700 505152 4752
rect 131028 4632 131080 4684
rect 219716 4632 219768 4684
rect 226340 4632 226392 4684
rect 299480 4632 299532 4684
rect 299572 4632 299624 4684
rect 320824 4632 320876 4684
rect 357348 4632 357400 4684
rect 442724 4632 442776 4684
rect 284300 4564 284352 4616
rect 326344 4564 326396 4616
rect 41052 4088 41104 4140
rect 183100 4088 183152 4140
rect 262956 4088 263008 4140
rect 487160 4088 487212 4140
rect 539508 4088 539560 4140
rect 575756 4088 575808 4140
rect 40684 4020 40736 4072
rect 189724 4020 189776 4072
rect 206284 4020 206336 4072
rect 219440 4020 219492 4072
rect 223028 4020 223080 4072
rect 234620 4020 234672 4072
rect 255228 4020 255280 4072
rect 492588 4020 492640 4072
rect 532608 4020 532660 4072
rect 542268 4020 542320 4072
rect 579068 4020 579120 4072
rect 40224 3952 40276 4004
rect 236276 3952 236328 4004
rect 276204 3952 276256 4004
rect 277308 3952 277360 4004
rect 286140 3952 286192 4004
rect 542544 3952 542596 4004
rect 547420 3952 547472 4004
rect 580172 3952 580224 4004
rect 38568 3884 38620 3936
rect 252836 3884 252888 3936
rect 272892 3884 272944 3936
rect 277400 3884 277452 3936
rect 279516 3884 279568 3936
rect 543096 3884 543148 3936
rect 40776 3816 40828 3868
rect 319444 3816 319496 3868
rect 324228 3816 324280 3868
rect 326068 3816 326120 3868
rect 400128 3816 400180 3868
rect 582380 3816 582432 3868
rect 38016 3748 38068 3800
rect 46572 3748 46624 3800
rect 59820 3748 59872 3800
rect 340880 3748 340932 3800
rect 367744 3748 367796 3800
rect 559196 3748 559248 3800
rect 39120 3680 39172 3732
rect 322756 3680 322808 3732
rect 326988 3680 327040 3732
rect 329564 3680 329616 3732
rect 332876 3680 332928 3732
rect 333888 3680 333940 3732
rect 336188 3680 336240 3732
rect 543188 3680 543240 3732
rect 3332 3612 3384 3664
rect 99380 3612 99432 3664
rect 113180 3612 113232 3664
rect 140780 3612 140832 3664
rect 146484 3612 146536 3664
rect 477500 3612 477552 3664
rect 505836 3612 505888 3664
rect 542636 3612 542688 3664
rect 41236 3544 41288 3596
rect 153108 3544 153160 3596
rect 156420 3544 156472 3596
rect 543556 3544 543608 3596
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 13268 3476 13320 3528
rect 13728 3476 13780 3528
rect 16580 3476 16632 3528
rect 17868 3476 17920 3528
rect 19892 3476 19944 3528
rect 20628 3476 20680 3528
rect 33140 3476 33192 3528
rect 34428 3476 34480 3528
rect 36636 3476 36688 3528
rect 37096 3476 37148 3528
rect 43260 3476 43312 3528
rect 44088 3476 44140 3528
rect 40500 3408 40552 3460
rect 469220 3476 469272 3528
rect 495900 3476 495952 3528
rect 545396 3476 545448 3528
rect 551284 3476 551336 3528
rect 552572 3476 552624 3528
rect 552664 3476 552716 3528
rect 569132 3476 569184 3528
rect 522580 3408 522632 3460
rect 535828 3408 535880 3460
rect 536748 3408 536800 3460
rect 572444 3408 572496 3460
rect 40960 3340 41012 3392
rect 166356 3340 166408 3392
rect 179604 3340 179656 3392
rect 198740 3340 198792 3392
rect 263508 3340 263560 3392
rect 485964 3340 486016 3392
rect 527088 3340 527140 3392
rect 562508 3340 562560 3392
rect 38476 3272 38528 3324
rect 40408 3204 40460 3256
rect 159732 3272 159784 3324
rect 149796 3204 149848 3256
rect 159364 3204 159416 3256
rect 289452 3272 289504 3324
rect 292948 3272 293000 3324
rect 295432 3272 295484 3324
rect 312820 3272 312872 3324
rect 517520 3272 517572 3324
rect 525892 3272 525944 3324
rect 543004 3272 543056 3324
rect 186412 3204 186464 3256
rect 187608 3204 187660 3256
rect 20 3136 72 3188
rect 1308 3136 1360 3188
rect 40868 3136 40920 3188
rect 133052 3136 133104 3188
rect 176292 3136 176344 3188
rect 41696 3068 41748 3120
rect 103060 3068 103112 3120
rect 131764 3068 131816 3120
rect 163044 3068 163096 3120
rect 182824 3068 182876 3120
rect 342812 3204 342864 3256
rect 360108 3204 360160 3256
rect 366180 3204 366232 3256
rect 402888 3204 402940 3256
rect 465908 3204 465960 3256
rect 532516 3204 532568 3256
rect 545212 3204 545264 3256
rect 193220 3136 193272 3188
rect 202788 3136 202840 3188
rect 346124 3136 346176 3188
rect 415308 3136 415360 3188
rect 429292 3136 429344 3188
rect 439504 3136 439556 3188
rect 446036 3136 446088 3188
rect 449348 3136 449400 3188
rect 449808 3136 449860 3188
rect 451924 3136 451976 3188
rect 455972 3136 456024 3188
rect 462596 3136 462648 3188
rect 523040 3136 523092 3188
rect 23204 3000 23256 3052
rect 64880 3000 64932 3052
rect 76564 3000 76616 3052
rect 131856 3000 131908 3052
rect 184848 3000 184900 3052
rect 306196 3068 306248 3120
rect 311808 3068 311860 3120
rect 399300 3068 399352 3120
rect 443644 3068 443696 3120
rect 502524 3068 502576 3120
rect 199660 3000 199712 3052
rect 284300 3000 284352 3052
rect 301504 3000 301556 3052
rect 416044 3000 416096 3052
rect 448428 3000 448480 3052
rect 472532 3000 472584 3052
rect 512644 3000 512696 3052
rect 513288 3000 513340 3052
rect 39948 2932 40000 2984
rect 77300 2932 77352 2984
rect 89812 2932 89864 2984
rect 120080 2932 120132 2984
rect 123116 2932 123168 2984
rect 147680 2932 147732 2984
rect 213828 2932 213880 2984
rect 216220 2932 216272 2984
rect 29828 2864 29880 2916
rect 62120 2864 62172 2916
rect 63132 2864 63184 2916
rect 92572 2864 92624 2916
rect 38660 2796 38712 2848
rect 53196 2796 53248 2848
rect 86960 2796 87012 2848
<< metal2 >>
rect 3118 703520 3230 704960
rect 3422 703760 3478 703769
rect 3422 703695 3478 703704
rect 3160 699786 3188 703520
rect 3436 702506 3464 703695
rect 6430 703520 6542 704960
rect 9742 703520 9854 704960
rect 13054 703520 13166 704960
rect 16366 703520 16478 704960
rect 19678 703520 19790 704960
rect 22990 703520 23102 704960
rect 26302 703520 26414 704960
rect 29614 703520 29726 704960
rect 32926 703520 33038 704960
rect 36422 703520 36534 704960
rect 39734 703520 39846 704960
rect 43046 703520 43158 704960
rect 46358 703520 46470 704960
rect 49670 703520 49782 704960
rect 52982 703520 53094 704960
rect 56294 703520 56406 704960
rect 59606 703520 59718 704960
rect 62918 703520 63030 704960
rect 66230 703520 66342 704960
rect 69542 703520 69654 704960
rect 73038 703520 73150 704960
rect 76350 703520 76462 704960
rect 79662 703520 79774 704960
rect 82974 703520 83086 704960
rect 86286 703520 86398 704960
rect 89598 703520 89710 704960
rect 92910 703520 93022 704960
rect 95252 703582 96108 703610
rect 3424 702500 3476 702506
rect 3424 702442 3476 702448
rect 6472 702434 6500 703520
rect 7748 702500 7800 702506
rect 7748 702442 7800 702448
rect 6472 702406 6868 702434
rect 3148 699780 3200 699786
rect 3148 699722 3200 699728
rect 6184 699780 6236 699786
rect 6184 699722 6236 699728
rect 3238 698592 3294 698601
rect 3238 698527 3294 698536
rect 3252 698358 3280 698527
rect 3240 698352 3292 698358
rect 3240 698294 3292 698300
rect 3146 693696 3202 693705
rect 3146 693631 3202 693640
rect 3160 692850 3188 693631
rect 3148 692844 3200 692850
rect 3148 692786 3200 692792
rect 3514 688800 3570 688809
rect 3514 688735 3570 688744
rect 3422 683904 3478 683913
rect 3422 683839 3478 683848
rect 3436 664630 3464 683839
rect 3424 664624 3476 664630
rect 3424 664566 3476 664572
rect 3422 664320 3478 664329
rect 3422 664255 3478 664264
rect 3436 663950 3464 664255
rect 3424 663944 3476 663950
rect 3424 663886 3476 663892
rect 3240 661632 3292 661638
rect 3240 661574 3292 661580
rect 3252 654294 3280 661574
rect 3332 659728 3384 659734
rect 3332 659670 3384 659676
rect 3240 654288 3292 654294
rect 3240 654230 3292 654236
rect 3344 649641 3372 659670
rect 3422 659424 3478 659433
rect 3422 659359 3478 659368
rect 3436 658442 3464 659359
rect 3424 658436 3476 658442
rect 3424 658378 3476 658384
rect 3422 654528 3478 654537
rect 3422 654463 3424 654472
rect 3476 654463 3478 654472
rect 3424 654434 3476 654440
rect 3424 654356 3476 654362
rect 3424 654298 3476 654304
rect 3330 649632 3386 649641
rect 3330 649567 3386 649576
rect 2780 640280 2832 640286
rect 2780 640222 2832 640228
rect 2792 639577 2820 640222
rect 2778 639568 2834 639577
rect 2778 639503 2834 639512
rect 2778 634672 2834 634681
rect 2778 634607 2834 634616
rect 2792 633554 2820 634607
rect 2780 633548 2832 633554
rect 2780 633490 2832 633496
rect 3332 615460 3384 615466
rect 3332 615402 3384 615408
rect 3344 615097 3372 615402
rect 3330 615088 3386 615097
rect 3330 615023 3386 615032
rect 3330 610192 3386 610201
rect 3330 610127 3332 610136
rect 3384 610127 3386 610136
rect 3332 610098 3384 610104
rect 3330 605296 3386 605305
rect 3330 605231 3386 605240
rect 3344 604518 3372 605231
rect 3332 604512 3384 604518
rect 3332 604454 3384 604460
rect 2780 601384 2832 601390
rect 2780 601326 2832 601332
rect 2792 600409 2820 601326
rect 2778 600400 2834 600409
rect 2778 600335 2834 600344
rect 3330 595504 3386 595513
rect 3330 595439 3386 595448
rect 3344 595066 3372 595439
rect 3332 595060 3384 595066
rect 3332 595002 3384 595008
rect 3332 593428 3384 593434
rect 3332 593370 3384 593376
rect 3148 590368 3200 590374
rect 3146 590336 3148 590345
rect 3200 590336 3202 590345
rect 3146 590271 3202 590280
rect 2780 585812 2832 585818
rect 2780 585754 2832 585760
rect 2792 585449 2820 585754
rect 2778 585440 2834 585449
rect 2778 585375 2834 585384
rect 3240 585200 3292 585206
rect 3240 585142 3292 585148
rect 3252 580553 3280 585142
rect 3238 580544 3294 580553
rect 3238 580479 3294 580488
rect 3240 578740 3292 578746
rect 3240 578682 3292 578688
rect 3146 575648 3202 575657
rect 3146 575583 3202 575592
rect 3054 570752 3110 570761
rect 3054 570687 3110 570696
rect 3068 570314 3096 570687
rect 3056 570308 3108 570314
rect 3056 570250 3108 570256
rect 2780 566024 2832 566030
rect 2780 565966 2832 565972
rect 2792 565865 2820 565966
rect 3056 565888 3108 565894
rect 2778 565856 2834 565865
rect 3056 565830 3108 565836
rect 2778 565791 2834 565800
rect 3068 547874 3096 565830
rect 3160 561678 3188 575583
rect 3148 561672 3200 561678
rect 3148 561614 3200 561620
rect 3146 560960 3202 560969
rect 3146 560895 3202 560904
rect 3160 560318 3188 560895
rect 3148 560312 3200 560318
rect 3148 560254 3200 560260
rect 3148 556164 3200 556170
rect 3148 556106 3200 556112
rect 3160 556073 3188 556106
rect 3146 556064 3202 556073
rect 3146 555999 3202 556008
rect 3146 551168 3202 551177
rect 3146 551103 3202 551112
rect 3160 550798 3188 551103
rect 3148 550792 3200 550798
rect 3148 550734 3200 550740
rect 3068 547846 3188 547874
rect 3160 546281 3188 547846
rect 3146 546272 3202 546281
rect 3146 546207 3202 546216
rect 3146 541376 3202 541385
rect 3146 541311 3202 541320
rect 3160 541006 3188 541311
rect 3148 541000 3200 541006
rect 3148 540942 3200 540948
rect 2778 531312 2834 531321
rect 2778 531247 2780 531256
rect 2832 531247 2834 531256
rect 2780 531218 2832 531224
rect 3146 521520 3202 521529
rect 3146 521455 3202 521464
rect 3160 520334 3188 521455
rect 3148 520328 3200 520334
rect 3148 520270 3200 520276
rect 3148 516724 3200 516730
rect 3148 516666 3200 516672
rect 3160 511737 3188 516666
rect 3146 511728 3202 511737
rect 3146 511663 3202 511672
rect 3146 487248 3202 487257
rect 3146 487183 3202 487192
rect 3054 482080 3110 482089
rect 3054 482015 3110 482024
rect 2962 477184 3018 477193
rect 2962 477119 3018 477128
rect 2976 471918 3004 477119
rect 2964 471912 3016 471918
rect 2964 471854 3016 471860
rect 3068 470594 3096 482015
rect 2976 470566 3096 470594
rect 2976 463690 3004 470566
rect 3160 467514 3188 487183
rect 3068 467486 3188 467514
rect 2964 463684 3016 463690
rect 2964 463626 3016 463632
rect 3068 459542 3096 467486
rect 3146 467392 3202 467401
rect 3146 467327 3148 467336
rect 3200 467327 3202 467336
rect 3148 467298 3200 467304
rect 3146 462496 3202 462505
rect 3146 462431 3148 462440
rect 3200 462431 3202 462440
rect 3148 462402 3200 462408
rect 3056 459536 3108 459542
rect 3056 459478 3108 459484
rect 3252 457609 3280 578682
rect 3238 457600 3294 457609
rect 3238 457535 3294 457544
rect 3240 452940 3292 452946
rect 3240 452882 3292 452888
rect 3252 452713 3280 452882
rect 3238 452704 3294 452713
rect 3238 452639 3294 452648
rect 3146 447808 3202 447817
rect 3146 447743 3202 447752
rect 3160 447166 3188 447743
rect 3148 447160 3200 447166
rect 3148 447102 3200 447108
rect 3240 444440 3292 444446
rect 3240 444382 3292 444388
rect 3252 442921 3280 444382
rect 3238 442912 3294 442921
rect 3238 442847 3294 442856
rect 3240 438864 3292 438870
rect 3240 438806 3292 438812
rect 3252 438025 3280 438806
rect 3238 438016 3294 438025
rect 3238 437951 3294 437960
rect 2962 433120 3018 433129
rect 2962 433055 3018 433064
rect 2976 431934 3004 433055
rect 2964 431928 3016 431934
rect 2964 431870 3016 431876
rect 3240 429072 3292 429078
rect 3240 429014 3292 429020
rect 3252 427961 3280 429014
rect 3238 427952 3294 427961
rect 3238 427887 3294 427896
rect 3240 423360 3292 423366
rect 3240 423302 3292 423308
rect 3252 423065 3280 423302
rect 3238 423056 3294 423065
rect 3238 422991 3294 423000
rect 3238 418160 3294 418169
rect 3238 418095 3240 418104
rect 3292 418095 3294 418104
rect 3240 418066 3292 418072
rect 3148 413704 3200 413710
rect 3148 413646 3200 413652
rect 3160 413273 3188 413646
rect 3146 413264 3202 413273
rect 3146 413199 3202 413208
rect 2780 408400 2832 408406
rect 2778 408368 2780 408377
rect 2832 408368 2834 408377
rect 2778 408303 2834 408312
rect 3240 404320 3292 404326
rect 3240 404262 3292 404268
rect 3252 403481 3280 404262
rect 3238 403472 3294 403481
rect 3238 403407 3294 403416
rect 3240 398608 3292 398614
rect 3238 398576 3240 398585
rect 3292 398576 3294 398585
rect 3238 398511 3294 398520
rect 2778 393680 2834 393689
rect 2778 393615 2780 393624
rect 2832 393615 2834 393624
rect 2780 393586 2832 393592
rect 2780 384804 2832 384810
rect 2780 384746 2832 384752
rect 2792 383897 2820 384746
rect 2778 383888 2834 383897
rect 2778 383823 2834 383832
rect 3238 368928 3294 368937
rect 3238 368863 3294 368872
rect 3252 368558 3280 368863
rect 3240 368552 3292 368558
rect 3240 368494 3292 368500
rect 3344 364041 3372 593370
rect 3330 364032 3386 364041
rect 3330 363967 3386 363976
rect 3148 354680 3200 354686
rect 3148 354622 3200 354628
rect 3160 354249 3188 354622
rect 3146 354240 3202 354249
rect 3146 354175 3202 354184
rect 2778 349344 2834 349353
rect 2778 349279 2834 349288
rect 2792 349246 2820 349279
rect 2780 349240 2832 349246
rect 2780 349182 2832 349188
rect 3330 344448 3386 344457
rect 3330 344383 3332 344392
rect 3384 344383 3386 344392
rect 3332 344354 3384 344360
rect 3330 339552 3386 339561
rect 3330 339487 3332 339496
rect 3384 339487 3386 339496
rect 3332 339458 3384 339464
rect 2964 334892 3016 334898
rect 2964 334834 3016 334840
rect 2976 334665 3004 334834
rect 2962 334656 3018 334665
rect 2962 334591 3018 334600
rect 3332 332648 3384 332654
rect 3332 332590 3384 332596
rect 3238 329760 3294 329769
rect 3238 329695 3294 329704
rect 3252 328778 3280 329695
rect 3240 328772 3292 328778
rect 3240 328714 3292 328720
rect 3344 319705 3372 332590
rect 3330 319696 3386 319705
rect 3330 319631 3386 319640
rect 3332 315988 3384 315994
rect 3332 315930 3384 315936
rect 3344 314809 3372 315930
rect 3330 314800 3386 314809
rect 3330 314735 3386 314744
rect 2964 314696 3016 314702
rect 2964 314638 3016 314644
rect 2976 309913 3004 314638
rect 3332 310548 3384 310554
rect 3332 310490 3384 310496
rect 2962 309904 3018 309913
rect 2962 309839 3018 309848
rect 2780 305040 2832 305046
rect 2778 305008 2780 305017
rect 2832 305008 2834 305017
rect 2778 304943 2834 304952
rect 3344 300121 3372 310490
rect 3330 300112 3386 300121
rect 3330 300047 3386 300056
rect 3332 295316 3384 295322
rect 3332 295258 3384 295264
rect 3344 295225 3372 295258
rect 3330 295216 3386 295225
rect 3330 295151 3386 295160
rect 3146 290320 3202 290329
rect 3146 290255 3202 290264
rect 3160 289882 3188 290255
rect 3148 289876 3200 289882
rect 3148 289818 3200 289824
rect 3238 285424 3294 285433
rect 3238 285359 3294 285368
rect 3148 266144 3200 266150
rect 3148 266086 3200 266092
rect 3160 265577 3188 266086
rect 3146 265568 3202 265577
rect 3146 265503 3202 265512
rect 3146 260672 3202 260681
rect 3146 260607 3202 260616
rect 3160 260234 3188 260607
rect 3148 260228 3200 260234
rect 3148 260170 3200 260176
rect 3146 226400 3202 226409
rect 3146 226335 3148 226344
rect 3200 226335 3202 226344
rect 3148 226306 3200 226312
rect 3148 220856 3200 220862
rect 3148 220798 3200 220804
rect 3054 216608 3110 216617
rect 3054 216543 3110 216552
rect 3068 211342 3096 216543
rect 3056 211336 3108 211342
rect 3056 211278 3108 211284
rect 3160 201657 3188 220798
rect 3146 201648 3202 201657
rect 3146 201583 3202 201592
rect 3146 196752 3202 196761
rect 3146 196687 3148 196696
rect 3200 196687 3202 196696
rect 3148 196658 3200 196664
rect 3146 186960 3202 186969
rect 3146 186895 3202 186904
rect 3160 186658 3188 186895
rect 3148 186652 3200 186658
rect 3148 186594 3200 186600
rect 3056 184952 3108 184958
rect 3056 184894 3108 184900
rect 3068 180794 3096 184894
rect 3148 182164 3200 182170
rect 3148 182106 3200 182112
rect 3160 182073 3188 182106
rect 3146 182064 3202 182073
rect 3146 181999 3202 182008
rect 3068 180766 3188 180794
rect 3054 177168 3110 177177
rect 3054 177103 3110 177112
rect 3068 177002 3096 177103
rect 3056 176996 3108 177002
rect 3056 176938 3108 176944
rect 3054 172272 3110 172281
rect 3054 172207 3110 172216
rect 3068 172174 3096 172207
rect 3056 172168 3108 172174
rect 3056 172110 3108 172116
rect 3160 167385 3188 180766
rect 3146 167376 3202 167385
rect 3146 167311 3202 167320
rect 2780 162512 2832 162518
rect 2778 162480 2780 162489
rect 2832 162480 2834 162489
rect 2778 162415 2834 162424
rect 2778 142624 2834 142633
rect 2778 142559 2834 142568
rect 2792 142390 2820 142559
rect 2780 142384 2832 142390
rect 2780 142326 2832 142332
rect 3252 132494 3280 285359
rect 3330 280528 3386 280537
rect 3330 280463 3332 280472
rect 3384 280463 3386 280472
rect 3332 280434 3384 280440
rect 3330 275632 3386 275641
rect 3330 275567 3386 275576
rect 3344 274718 3372 275567
rect 3332 274712 3384 274718
rect 3332 274654 3384 274660
rect 3330 270736 3386 270745
rect 3330 270671 3386 270680
rect 3160 132466 3280 132494
rect 3160 125662 3188 132466
rect 3240 128308 3292 128314
rect 3240 128250 3292 128256
rect 3252 127945 3280 128250
rect 3238 127936 3294 127945
rect 3238 127871 3294 127880
rect 3148 125656 3200 125662
rect 3148 125598 3200 125604
rect 3054 113248 3110 113257
rect 3054 113183 3056 113192
rect 3108 113183 3110 113192
rect 3056 113154 3108 113160
rect 3344 109614 3372 270671
rect 3436 157321 3464 654298
rect 3528 651370 3556 688735
rect 3882 679008 3938 679017
rect 3882 678943 3938 678952
rect 3698 674112 3754 674121
rect 3698 674047 3754 674056
rect 3608 661156 3660 661162
rect 3608 661098 3660 661104
rect 3620 654430 3648 661098
rect 3608 654424 3660 654430
rect 3608 654366 3660 654372
rect 3608 654288 3660 654294
rect 3608 654230 3660 654236
rect 3516 651364 3568 651370
rect 3516 651306 3568 651312
rect 3516 630624 3568 630630
rect 3516 630566 3568 630572
rect 3528 629785 3556 630566
rect 3514 629776 3570 629785
rect 3514 629711 3570 629720
rect 3516 618248 3568 618254
rect 3516 618190 3568 618196
rect 3528 507362 3556 618190
rect 3620 507482 3648 654230
rect 3712 647222 3740 674047
rect 3790 669216 3846 669225
rect 3790 669151 3846 669160
rect 3700 647216 3752 647222
rect 3700 647158 3752 647164
rect 3698 644464 3754 644473
rect 3698 644399 3754 644408
rect 3712 601662 3740 644399
rect 3804 643074 3832 669151
rect 3896 660346 3924 678943
rect 5172 665100 5224 665106
rect 5172 665042 5224 665048
rect 5080 664828 5132 664834
rect 5080 664770 5132 664776
rect 4988 664216 5040 664222
rect 4988 664158 5040 664164
rect 4804 664080 4856 664086
rect 4804 664022 4856 664028
rect 4712 663876 4764 663882
rect 4712 663818 4764 663824
rect 4068 661768 4120 661774
rect 4068 661710 4120 661716
rect 3976 661496 4028 661502
rect 3976 661438 4028 661444
rect 3884 660340 3936 660346
rect 3884 660282 3936 660288
rect 3792 643068 3844 643074
rect 3792 643010 3844 643016
rect 3882 624880 3938 624889
rect 3882 624815 3938 624824
rect 3792 619540 3844 619546
rect 3792 619482 3844 619488
rect 3700 601656 3752 601662
rect 3700 601598 3752 601604
rect 3700 579692 3752 579698
rect 3700 579634 3752 579640
rect 3712 516730 3740 579634
rect 3700 516724 3752 516730
rect 3700 516666 3752 516672
rect 3698 516624 3754 516633
rect 3698 516559 3754 516568
rect 3712 516458 3740 516559
rect 3700 516452 3752 516458
rect 3700 516394 3752 516400
rect 3608 507476 3660 507482
rect 3608 507418 3660 507424
rect 3528 507334 3740 507362
rect 3608 507272 3660 507278
rect 3608 507214 3660 507220
rect 3516 507204 3568 507210
rect 3516 507146 3568 507152
rect 3528 506841 3556 507146
rect 3514 506832 3570 506841
rect 3514 506767 3570 506776
rect 3514 492144 3570 492153
rect 3514 492079 3570 492088
rect 3528 485790 3556 492079
rect 3516 485784 3568 485790
rect 3516 485726 3568 485732
rect 3514 472288 3570 472297
rect 3514 472223 3570 472232
rect 3528 472054 3556 472223
rect 3516 472048 3568 472054
rect 3516 471990 3568 471996
rect 3516 471912 3568 471918
rect 3516 471854 3568 471860
rect 3422 157312 3478 157321
rect 3422 157247 3478 157256
rect 3424 147620 3476 147626
rect 3424 147562 3476 147568
rect 3436 147529 3464 147562
rect 3422 147520 3478 147529
rect 3422 147455 3478 147464
rect 3422 137728 3478 137737
rect 3422 137663 3478 137672
rect 3436 137562 3464 137663
rect 3424 137556 3476 137562
rect 3424 137498 3476 137504
rect 3422 132832 3478 132841
rect 3422 132767 3478 132776
rect 3332 109608 3384 109614
rect 3332 109550 3384 109556
rect 3148 108724 3200 108730
rect 3148 108666 3200 108672
rect 3160 108361 3188 108666
rect 3146 108352 3202 108361
rect 3146 108287 3202 108296
rect 3332 103488 3384 103494
rect 3332 103430 3384 103436
rect 3344 103193 3372 103430
rect 3330 103184 3386 103193
rect 3330 103119 3386 103128
rect 2778 93392 2834 93401
rect 2778 93327 2834 93336
rect 2792 92818 2820 93327
rect 2780 92812 2832 92818
rect 2780 92754 2832 92760
rect 3330 83600 3386 83609
rect 3330 83535 3386 83544
rect 3344 82890 3372 83535
rect 3332 82884 3384 82890
rect 3332 82826 3384 82832
rect 2780 78736 2832 78742
rect 2778 78704 2780 78713
rect 2832 78704 2834 78713
rect 2778 78639 2834 78648
rect 3332 74520 3384 74526
rect 3332 74462 3384 74468
rect 3344 73817 3372 74462
rect 3330 73808 3386 73817
rect 3330 73743 3386 73752
rect 3332 68944 3384 68950
rect 3330 68912 3332 68921
rect 3384 68912 3386 68921
rect 3330 68847 3386 68856
rect 2780 64048 2832 64054
rect 2778 64016 2780 64025
rect 2832 64016 2834 64025
rect 2778 63951 2834 63960
rect 3330 54224 3386 54233
rect 3330 54159 3386 54168
rect 2778 49056 2834 49065
rect 2778 48991 2834 49000
rect 2792 48346 2820 48991
rect 2780 48340 2832 48346
rect 2780 48282 2832 48288
rect 3240 44804 3292 44810
rect 3240 44746 3292 44752
rect 1308 39772 1360 39778
rect 1308 39714 1360 39720
rect 1320 3194 1348 39714
rect 2780 39704 2832 39710
rect 2780 39646 2832 39652
rect 2792 39273 2820 39646
rect 2778 39264 2834 39273
rect 2778 39199 2834 39208
rect 3252 39001 3280 44746
rect 3344 41410 3372 54159
rect 3332 41404 3384 41410
rect 3332 41346 3384 41352
rect 3436 40798 3464 132767
rect 3528 44810 3556 471854
rect 3620 255785 3648 507214
rect 3712 501945 3740 507334
rect 3698 501936 3754 501945
rect 3698 501871 3754 501880
rect 3698 497040 3754 497049
rect 3698 496975 3754 496984
rect 3606 255776 3662 255785
rect 3606 255711 3662 255720
rect 3608 246152 3660 246158
rect 3608 246094 3660 246100
rect 3620 245993 3648 246094
rect 3606 245984 3662 245993
rect 3606 245919 3662 245928
rect 3608 241120 3660 241126
rect 3606 241088 3608 241097
rect 3660 241088 3662 241097
rect 3606 241023 3662 241032
rect 3608 236224 3660 236230
rect 3606 236192 3608 236201
rect 3660 236192 3662 236201
rect 3606 236127 3662 236136
rect 3608 212492 3660 212498
rect 3608 212434 3660 212440
rect 3620 211449 3648 212434
rect 3606 211440 3662 211449
rect 3606 211375 3662 211384
rect 3608 211336 3660 211342
rect 3608 211278 3660 211284
rect 3620 139466 3648 211278
rect 3608 139460 3660 139466
rect 3608 139402 3660 139408
rect 3712 125594 3740 496975
rect 3804 250889 3832 619482
rect 3896 589286 3924 624815
rect 3884 589280 3936 589286
rect 3884 589222 3936 589228
rect 3884 564460 3936 564466
rect 3884 564402 3936 564408
rect 3790 250880 3846 250889
rect 3790 250815 3846 250824
rect 3896 231305 3924 564402
rect 3988 388793 4016 661438
rect 3974 388784 4030 388793
rect 3974 388719 4030 388728
rect 3974 373824 4030 373833
rect 3974 373759 4030 373768
rect 3882 231296 3938 231305
rect 3882 231231 3938 231240
rect 3882 221504 3938 221513
rect 3882 221439 3938 221448
rect 3790 206544 3846 206553
rect 3790 206479 3846 206488
rect 3804 153202 3832 206479
rect 3896 201482 3924 221439
rect 3884 201476 3936 201482
rect 3884 201418 3936 201424
rect 3882 191856 3938 191865
rect 3882 191791 3938 191800
rect 3896 172514 3924 191791
rect 3884 172508 3936 172514
rect 3884 172450 3936 172456
rect 3792 153196 3844 153202
rect 3792 153138 3844 153144
rect 3700 125588 3752 125594
rect 3700 125530 3752 125536
rect 3606 123040 3662 123049
rect 3606 122975 3608 122984
rect 3660 122975 3662 122984
rect 3608 122946 3660 122952
rect 3606 118144 3662 118153
rect 3606 118079 3662 118088
rect 3620 117366 3648 118079
rect 3608 117360 3660 117366
rect 3608 117302 3660 117308
rect 3606 88496 3662 88505
rect 3606 88431 3662 88440
rect 3516 44804 3568 44810
rect 3516 44746 3568 44752
rect 3620 44690 3648 88431
rect 3700 59424 3752 59430
rect 3700 59366 3752 59372
rect 3528 44662 3648 44690
rect 3424 40792 3476 40798
rect 3424 40734 3476 40740
rect 3528 39098 3556 44662
rect 3608 44532 3660 44538
rect 3608 44474 3660 44480
rect 3620 39846 3648 44474
rect 3608 39840 3660 39846
rect 3608 39782 3660 39788
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3238 38992 3294 39001
rect 3238 38927 3294 38936
rect 3424 34400 3476 34406
rect 3422 34368 3424 34377
rect 3476 34368 3478 34377
rect 3422 34303 3478 34312
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3252 24585 3280 24686
rect 3238 24576 3294 24585
rect 3238 24511 3294 24520
rect 3712 19689 3740 59366
rect 3790 59120 3846 59129
rect 3790 59055 3846 59064
rect 3804 44538 3832 59055
rect 3792 44532 3844 44538
rect 3792 44474 3844 44480
rect 3988 44418 4016 373759
rect 4080 359145 4108 661710
rect 4620 629944 4672 629950
rect 4620 629886 4672 629892
rect 4632 618254 4660 629886
rect 4620 618248 4672 618254
rect 4620 618190 4672 618196
rect 4724 601390 4752 663818
rect 4712 601384 4764 601390
rect 4712 601326 4764 601332
rect 4160 582344 4212 582350
rect 4160 582286 4212 582292
rect 4172 579698 4200 582286
rect 4252 580984 4304 580990
rect 4252 580926 4304 580932
rect 4160 579692 4212 579698
rect 4160 579634 4212 579640
rect 4264 578746 4292 580926
rect 4252 578740 4304 578746
rect 4252 578682 4304 578688
rect 4712 573776 4764 573782
rect 4712 573718 4764 573724
rect 4344 568540 4396 568546
rect 4344 568482 4396 568488
rect 4356 565894 4384 568482
rect 4344 565888 4396 565894
rect 4344 565830 4396 565836
rect 4724 564466 4752 573718
rect 4712 564460 4764 564466
rect 4712 564402 4764 564408
rect 4066 359136 4122 359145
rect 4066 359071 4122 359080
rect 4066 324864 4122 324873
rect 4066 324799 4122 324808
rect 3804 44390 4016 44418
rect 3804 40186 3832 44390
rect 4080 44282 4108 324799
rect 4712 125588 4764 125594
rect 4712 125530 4764 125536
rect 4724 118658 4752 125530
rect 4712 118652 4764 118658
rect 4712 118594 4764 118600
rect 4816 64054 4844 664022
rect 4896 661836 4948 661842
rect 4896 661778 4948 661784
rect 4908 640286 4936 661778
rect 4896 640280 4948 640286
rect 4896 640222 4948 640228
rect 4896 633548 4948 633554
rect 4896 633490 4948 633496
rect 4804 64048 4856 64054
rect 4804 63990 4856 63996
rect 4712 48340 4764 48346
rect 4712 48282 4764 48288
rect 3988 44254 4108 44282
rect 3882 43480 3938 43489
rect 3882 43415 3938 43424
rect 3792 40180 3844 40186
rect 3792 40122 3844 40128
rect 3896 29481 3924 43415
rect 3988 40390 4016 44254
rect 4066 44160 4122 44169
rect 4122 44118 4200 44146
rect 4066 44095 4122 44104
rect 4172 42294 4200 44118
rect 4160 42288 4212 42294
rect 4160 42230 4212 42236
rect 4724 40662 4752 48282
rect 4804 43444 4856 43450
rect 4804 43386 4856 43392
rect 4712 40656 4764 40662
rect 4712 40598 4764 40604
rect 3976 40384 4028 40390
rect 3976 40326 4028 40332
rect 3882 29472 3938 29481
rect 3882 29407 3938 29416
rect 3698 19680 3754 19689
rect 3698 19615 3754 19624
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3436 14793 3464 15098
rect 3422 14784 3478 14793
rect 3422 14719 3478 14728
rect 2964 9920 3016 9926
rect 2962 9888 2964 9897
rect 3016 9888 3018 9897
rect 2962 9823 3018 9832
rect 4816 5302 4844 43386
rect 4908 41002 4936 633490
rect 5000 585818 5028 664158
rect 4988 585812 5040 585818
rect 4988 585754 5040 585760
rect 4988 574116 5040 574122
rect 4988 574058 5040 574064
rect 4896 40996 4948 41002
rect 4896 40938 4948 40944
rect 5000 39710 5028 574058
rect 5092 162518 5120 664770
rect 5184 408406 5212 665042
rect 5264 663536 5316 663542
rect 5264 663478 5316 663484
rect 5172 408400 5224 408406
rect 5172 408342 5224 408348
rect 5172 393644 5224 393650
rect 5172 393586 5224 393592
rect 5080 162512 5132 162518
rect 5080 162454 5132 162460
rect 5080 142384 5132 142390
rect 5080 142326 5132 142332
rect 5092 40322 5120 142326
rect 5080 40316 5132 40322
rect 5080 40258 5132 40264
rect 5184 39914 5212 393586
rect 5276 384810 5304 663478
rect 5448 662924 5500 662930
rect 5448 662866 5500 662872
rect 5356 662856 5408 662862
rect 5356 662798 5408 662804
rect 5368 531282 5396 662798
rect 5460 566030 5488 662866
rect 5540 634772 5592 634778
rect 5540 634714 5592 634720
rect 5552 629950 5580 634714
rect 5540 629944 5592 629950
rect 5540 629886 5592 629892
rect 5540 597576 5592 597582
rect 5540 597518 5592 597524
rect 5552 593434 5580 597518
rect 5540 593428 5592 593434
rect 5540 593370 5592 593376
rect 5448 566024 5500 566030
rect 5448 565966 5500 565972
rect 5356 531276 5408 531282
rect 5356 531218 5408 531224
rect 5264 384804 5316 384810
rect 5264 384746 5316 384752
rect 5264 349240 5316 349246
rect 5264 349182 5316 349188
rect 5276 41070 5304 349182
rect 5356 346452 5408 346458
rect 5356 346394 5408 346400
rect 5368 305046 5396 346394
rect 5356 305040 5408 305046
rect 5356 304982 5408 304988
rect 5448 201476 5500 201482
rect 5448 201418 5500 201424
rect 5460 194546 5488 201418
rect 5448 194540 5500 194546
rect 5448 194482 5500 194488
rect 5448 172508 5500 172514
rect 5448 172450 5500 172456
rect 5460 165578 5488 172450
rect 5448 165572 5500 165578
rect 5448 165514 5500 165520
rect 5356 153196 5408 153202
rect 5356 153138 5408 153144
rect 5368 142154 5396 153138
rect 5368 142126 5580 142154
rect 5552 140350 5580 142126
rect 5540 140344 5592 140350
rect 5540 140286 5592 140292
rect 6092 139392 6144 139398
rect 6092 139334 6144 139340
rect 6104 131102 6132 139334
rect 6092 131096 6144 131102
rect 6092 131038 6144 131044
rect 5540 125588 5592 125594
rect 5540 125530 5592 125536
rect 5552 121038 5580 125530
rect 5540 121032 5592 121038
rect 5540 120974 5592 120980
rect 5540 118652 5592 118658
rect 5540 118594 5592 118600
rect 5552 115666 5580 118594
rect 5540 115660 5592 115666
rect 5540 115602 5592 115608
rect 6092 113212 6144 113218
rect 6092 113154 6144 113160
rect 5356 109608 5408 109614
rect 5356 109550 5408 109556
rect 5368 107642 5396 109550
rect 5356 107636 5408 107642
rect 5356 107578 5408 107584
rect 5356 92812 5408 92818
rect 5356 92754 5408 92760
rect 5264 41064 5316 41070
rect 5264 41006 5316 41012
rect 5368 40730 5396 92754
rect 5448 78736 5500 78742
rect 5448 78678 5500 78684
rect 5356 40724 5408 40730
rect 5356 40666 5408 40672
rect 5460 40254 5488 78678
rect 5448 40248 5500 40254
rect 5448 40190 5500 40196
rect 5172 39908 5224 39914
rect 5172 39850 5224 39856
rect 4988 39704 5040 39710
rect 4988 39646 5040 39652
rect 6104 39302 6132 113154
rect 6196 40361 6224 699722
rect 6552 664420 6604 664426
rect 6552 664362 6604 664368
rect 6368 661564 6420 661570
rect 6368 661506 6420 661512
rect 6274 661192 6330 661201
rect 6274 661127 6330 661136
rect 6182 40352 6238 40361
rect 6182 40287 6238 40296
rect 6092 39296 6144 39302
rect 6092 39238 6144 39244
rect 6288 9926 6316 661127
rect 6380 24750 6408 661506
rect 6460 659864 6512 659870
rect 6460 659806 6512 659812
rect 6472 334898 6500 659806
rect 6564 590374 6592 664362
rect 6644 661972 6696 661978
rect 6644 661914 6696 661920
rect 6552 590368 6604 590374
rect 6552 590310 6604 590316
rect 6552 550792 6604 550798
rect 6552 550734 6604 550740
rect 6460 334892 6512 334898
rect 6460 334834 6512 334840
rect 6460 328772 6512 328778
rect 6460 328714 6512 328720
rect 6472 38826 6500 328714
rect 6564 270502 6592 550734
rect 6656 413710 6684 661914
rect 6840 661026 6868 702406
rect 7656 664148 7708 664154
rect 7656 664090 7708 664096
rect 6828 661020 6880 661026
rect 6828 660962 6880 660968
rect 6736 658436 6788 658442
rect 6736 658378 6788 658384
rect 6748 597514 6776 658378
rect 7564 654492 7616 654498
rect 7564 654434 7616 654440
rect 6736 597508 6788 597514
rect 6736 597450 6788 597456
rect 6736 529984 6788 529990
rect 6736 529926 6788 529932
rect 6748 429078 6776 529926
rect 6736 429072 6788 429078
rect 6736 429014 6788 429020
rect 6644 413704 6696 413710
rect 6644 413646 6696 413652
rect 6828 398880 6880 398886
rect 6828 398822 6880 398828
rect 6644 350600 6696 350606
rect 6644 350542 6696 350548
rect 6552 270496 6604 270502
rect 6552 270438 6604 270444
rect 6552 226364 6604 226370
rect 6552 226306 6604 226312
rect 6564 40866 6592 226306
rect 6656 108730 6684 350542
rect 6736 176996 6788 177002
rect 6736 176938 6788 176944
rect 6644 108724 6696 108730
rect 6644 108666 6696 108672
rect 6644 107636 6696 107642
rect 6644 107578 6696 107584
rect 6656 102678 6684 107578
rect 6644 102672 6696 102678
rect 6644 102614 6696 102620
rect 6552 40860 6604 40866
rect 6552 40802 6604 40808
rect 6748 40118 6776 176938
rect 6736 40112 6788 40118
rect 6736 40054 6788 40060
rect 6460 38820 6512 38826
rect 6460 38762 6512 38768
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6840 6914 6868 398822
rect 7472 121032 7524 121038
rect 7472 120974 7524 120980
rect 7484 117094 7512 120974
rect 7472 117088 7524 117094
rect 7472 117030 7524 117036
rect 7472 115660 7524 115666
rect 7472 115602 7524 115608
rect 7484 109682 7512 115602
rect 7472 109676 7524 109682
rect 7472 109618 7524 109624
rect 7472 102672 7524 102678
rect 7472 102614 7524 102620
rect 7484 99074 7512 102614
rect 7472 99068 7524 99074
rect 7472 99010 7524 99016
rect 7576 41274 7604 654434
rect 7668 630630 7696 664090
rect 7656 630624 7708 630630
rect 7656 630566 7708 630572
rect 7656 600296 7708 600302
rect 7656 600238 7708 600244
rect 7668 581058 7696 600238
rect 7656 581052 7708 581058
rect 7656 580994 7708 581000
rect 7656 570308 7708 570314
rect 7656 570250 7708 570256
rect 7564 41268 7616 41274
rect 7564 41210 7616 41216
rect 7668 38690 7696 570250
rect 7760 539578 7788 702442
rect 9784 700126 9812 703520
rect 16408 702434 16436 703520
rect 16408 702406 16528 702434
rect 9772 700120 9824 700126
rect 9772 700062 9824 700068
rect 10968 700120 11020 700126
rect 10968 700062 11020 700068
rect 10324 692844 10376 692850
rect 10324 692786 10376 692792
rect 7932 664896 7984 664902
rect 7932 664838 7984 664844
rect 8942 664864 8998 664873
rect 7840 662040 7892 662046
rect 7840 661982 7892 661988
rect 7748 539572 7800 539578
rect 7748 539514 7800 539520
rect 7748 467356 7800 467362
rect 7748 467298 7800 467304
rect 7760 40934 7788 467298
rect 7852 236230 7880 661982
rect 7944 507210 7972 664838
rect 8942 664799 8998 664808
rect 8116 662108 8168 662114
rect 8116 662050 8168 662056
rect 8024 590640 8076 590646
rect 8024 590582 8076 590588
rect 8036 582418 8064 590582
rect 8024 582412 8076 582418
rect 8024 582354 8076 582360
rect 8024 574184 8076 574190
rect 8024 574126 8076 574132
rect 8036 568614 8064 574126
rect 8024 568608 8076 568614
rect 8024 568550 8076 568556
rect 7932 507204 7984 507210
rect 7932 507146 7984 507152
rect 8024 488572 8076 488578
rect 8024 488514 8076 488520
rect 7932 462460 7984 462466
rect 7932 462402 7984 462408
rect 7840 236224 7892 236230
rect 7840 236166 7892 236172
rect 7840 186652 7892 186658
rect 7840 186594 7892 186600
rect 7852 41342 7880 186594
rect 7840 41336 7892 41342
rect 7840 41278 7892 41284
rect 7748 40928 7800 40934
rect 7748 40870 7800 40876
rect 7944 40458 7972 462402
rect 8036 68950 8064 488514
rect 8128 246158 8156 662050
rect 8484 637560 8536 637566
rect 8484 637502 8536 637508
rect 8496 634846 8524 637502
rect 8484 634840 8536 634846
rect 8484 634782 8536 634788
rect 8208 622396 8260 622402
rect 8208 622338 8260 622344
rect 8220 619546 8248 622338
rect 8208 619540 8260 619546
rect 8208 619482 8260 619488
rect 8852 610156 8904 610162
rect 8852 610098 8904 610104
rect 8208 604580 8260 604586
rect 8208 604522 8260 604528
rect 8220 597582 8248 604522
rect 8208 597576 8260 597582
rect 8208 597518 8260 597524
rect 8300 591116 8352 591122
rect 8300 591058 8352 591064
rect 8312 590594 8340 591058
rect 8220 590566 8340 590594
rect 8220 585206 8248 590566
rect 8208 585200 8260 585206
rect 8208 585142 8260 585148
rect 8300 577176 8352 577182
rect 8300 577118 8352 577124
rect 8312 573782 8340 577118
rect 8300 573776 8352 573782
rect 8300 573718 8352 573724
rect 8864 499526 8892 610098
rect 8852 499520 8904 499526
rect 8852 499462 8904 499468
rect 8116 246152 8168 246158
rect 8116 246094 8168 246100
rect 8116 194540 8168 194546
rect 8116 194482 8168 194488
rect 8128 173874 8156 194482
rect 8116 173868 8168 173874
rect 8116 173810 8168 173816
rect 8116 165572 8168 165578
rect 8116 165514 8168 165520
rect 8128 144906 8156 165514
rect 8116 144900 8168 144906
rect 8116 144842 8168 144848
rect 8208 140344 8260 140350
rect 8208 140286 8260 140292
rect 8220 137902 8248 140286
rect 8208 137896 8260 137902
rect 8208 137838 8260 137844
rect 8116 137556 8168 137562
rect 8116 137498 8168 137504
rect 8024 68944 8076 68950
rect 8024 68886 8076 68892
rect 7932 40452 7984 40458
rect 7932 40394 7984 40400
rect 8128 39438 8156 137498
rect 8852 131096 8904 131102
rect 8852 131038 8904 131044
rect 8864 126954 8892 131038
rect 8852 126948 8904 126954
rect 8852 126890 8904 126896
rect 8208 123004 8260 123010
rect 8208 122946 8260 122952
rect 8220 39574 8248 122946
rect 8852 99068 8904 99074
rect 8852 99010 8904 99016
rect 8864 96626 8892 99010
rect 8852 96620 8904 96626
rect 8852 96562 8904 96568
rect 8208 39568 8260 39574
rect 8208 39510 8260 39516
rect 8116 39432 8168 39438
rect 8116 39374 8168 39380
rect 7656 38684 7708 38690
rect 7656 38626 7708 38632
rect 8956 34406 8984 664799
rect 9588 664692 9640 664698
rect 9588 664634 9640 664640
rect 9312 664488 9364 664494
rect 9312 664430 9364 664436
rect 9128 662584 9180 662590
rect 9128 662526 9180 662532
rect 9036 609952 9088 609958
rect 9036 609894 9088 609900
rect 9048 600302 9076 609894
rect 9036 600296 9088 600302
rect 9036 600238 9088 600244
rect 9036 583772 9088 583778
rect 9036 583714 9088 583720
rect 9048 574190 9076 583714
rect 9036 574184 9088 574190
rect 9036 574126 9088 574132
rect 9036 516452 9088 516458
rect 9036 516394 9088 516400
rect 9048 40594 9076 516394
rect 9140 241126 9168 662526
rect 9220 595060 9272 595066
rect 9220 595002 9272 595008
rect 9128 241120 9180 241126
rect 9128 241062 9180 241068
rect 9232 208350 9260 595002
rect 9324 398614 9352 664430
rect 9404 664284 9456 664290
rect 9404 664226 9456 664232
rect 9416 418130 9444 664226
rect 9496 662992 9548 662998
rect 9496 662934 9548 662940
rect 9508 423366 9536 662934
rect 9600 452946 9628 664634
rect 10232 594856 10284 594862
rect 10232 594798 10284 594804
rect 10244 591122 10272 594798
rect 10232 591116 10284 591122
rect 10232 591058 10284 591064
rect 9680 586492 9732 586498
rect 9680 586434 9732 586440
rect 9692 583778 9720 586434
rect 9680 583772 9732 583778
rect 9680 583714 9732 583720
rect 9588 452940 9640 452946
rect 9588 452882 9640 452888
rect 9496 423360 9548 423366
rect 9496 423302 9548 423308
rect 9404 418124 9456 418130
rect 9404 418066 9456 418072
rect 9588 412684 9640 412690
rect 9588 412626 9640 412632
rect 9312 398608 9364 398614
rect 9312 398550 9364 398556
rect 9312 344412 9364 344418
rect 9312 344354 9364 344360
rect 9220 208344 9272 208350
rect 9220 208286 9272 208292
rect 9128 196716 9180 196722
rect 9128 196658 9180 196664
rect 9140 41138 9168 196658
rect 9220 172168 9272 172174
rect 9220 172110 9272 172116
rect 9128 41132 9180 41138
rect 9128 41074 9180 41080
rect 9036 40588 9088 40594
rect 9036 40530 9088 40536
rect 9232 39642 9260 172110
rect 9220 39636 9272 39642
rect 9220 39578 9272 39584
rect 9324 39506 9352 344354
rect 9404 339516 9456 339522
rect 9404 339458 9456 339464
rect 9312 39500 9364 39506
rect 9312 39442 9364 39448
rect 9416 39234 9444 339458
rect 9496 280492 9548 280498
rect 9496 280434 9548 280440
rect 9508 39710 9536 280434
rect 9600 266150 9628 412626
rect 9588 266144 9640 266150
rect 9588 266086 9640 266092
rect 9588 260228 9640 260234
rect 9588 260170 9640 260176
rect 9600 168366 9628 260170
rect 9588 168360 9640 168366
rect 9588 168302 9640 168308
rect 9588 137896 9640 137902
rect 9588 137838 9640 137844
rect 9600 126886 9628 137838
rect 9588 126880 9640 126886
rect 9588 126822 9640 126828
rect 9588 117088 9640 117094
rect 9588 117030 9640 117036
rect 9600 110498 9628 117030
rect 9588 110492 9640 110498
rect 9588 110434 9640 110440
rect 10336 40225 10364 692786
rect 10600 664964 10652 664970
rect 10600 664906 10652 664912
rect 10416 664012 10468 664018
rect 10416 663954 10468 663960
rect 10428 74526 10456 663954
rect 10508 663944 10560 663950
rect 10508 663886 10560 663892
rect 10416 74520 10468 74526
rect 10416 74462 10468 74468
rect 10322 40216 10378 40225
rect 10322 40151 10378 40160
rect 10520 40089 10548 663886
rect 10612 128314 10640 664906
rect 10876 664556 10928 664562
rect 10876 664498 10928 664504
rect 10692 663944 10744 663950
rect 10692 663886 10744 663892
rect 10704 182170 10732 663886
rect 10784 596828 10836 596834
rect 10784 596770 10836 596776
rect 10796 577182 10824 596770
rect 10784 577176 10836 577182
rect 10784 577118 10836 577124
rect 10784 472048 10836 472054
rect 10784 471990 10836 471996
rect 10692 182164 10744 182170
rect 10692 182106 10744 182112
rect 10600 128308 10652 128314
rect 10600 128250 10652 128256
rect 10600 109676 10652 109682
rect 10600 109618 10652 109624
rect 10612 98870 10640 109618
rect 10796 109002 10824 471990
rect 10888 354686 10916 664498
rect 10980 660249 11008 700062
rect 11704 664352 11756 664358
rect 11704 664294 11756 664300
rect 10966 660240 11022 660249
rect 10966 660175 11022 660184
rect 11060 638988 11112 638994
rect 11060 638930 11112 638936
rect 11072 637634 11100 638930
rect 11060 637628 11112 637634
rect 11060 637570 11112 637576
rect 11336 608252 11388 608258
rect 11336 608194 11388 608200
rect 11348 604586 11376 608194
rect 11336 604580 11388 604586
rect 11336 604522 11388 604528
rect 11428 601792 11480 601798
rect 11428 601734 11480 601740
rect 10968 601724 11020 601730
rect 10968 601666 11020 601672
rect 10980 590714 11008 601666
rect 11440 596834 11468 601734
rect 11428 596828 11480 596834
rect 11428 596770 11480 596776
rect 10968 590708 11020 590714
rect 10968 590650 11020 590656
rect 11716 438870 11744 664294
rect 13820 645924 13872 645930
rect 13820 645866 13872 645872
rect 13832 644474 13860 645866
rect 13740 644446 13860 644474
rect 13740 638994 13768 644446
rect 13728 638988 13780 638994
rect 13728 638930 13780 638936
rect 15844 629672 15896 629678
rect 15844 629614 15896 629620
rect 15856 622470 15884 629614
rect 15844 622464 15896 622470
rect 15844 622406 15896 622412
rect 15844 619608 15896 619614
rect 15844 619550 15896 619556
rect 14464 619540 14516 619546
rect 14464 619482 14516 619488
rect 13820 614168 13872 614174
rect 13820 614110 13872 614116
rect 13832 611402 13860 614110
rect 13740 611374 13860 611402
rect 13740 608258 13768 611374
rect 13728 608252 13780 608258
rect 13728 608194 13780 608200
rect 13820 604648 13872 604654
rect 13820 604590 13872 604596
rect 13832 601730 13860 604590
rect 13912 604580 13964 604586
rect 13912 604522 13964 604528
rect 13924 601798 13952 604522
rect 13912 601792 13964 601798
rect 13912 601734 13964 601740
rect 13820 601724 13872 601730
rect 13820 601666 13872 601672
rect 13084 600296 13136 600302
rect 13084 600238 13136 600244
rect 13096 594862 13124 600238
rect 13084 594856 13136 594862
rect 13084 594798 13136 594804
rect 14476 586566 14504 619482
rect 15856 614174 15884 619550
rect 15844 614168 15896 614174
rect 15844 614110 15896 614116
rect 15844 611176 15896 611182
rect 15844 611118 15896 611124
rect 15200 605124 15252 605130
rect 15200 605066 15252 605072
rect 15212 600370 15240 605066
rect 15856 604586 15884 611118
rect 15844 604580 15896 604586
rect 15844 604522 15896 604528
rect 15200 600364 15252 600370
rect 15200 600306 15252 600312
rect 14464 586560 14516 586566
rect 14464 586502 14516 586508
rect 14464 560312 14516 560318
rect 14464 560254 14516 560260
rect 13084 447160 13136 447166
rect 13084 447102 13136 447108
rect 11704 438864 11756 438870
rect 11704 438806 11756 438812
rect 10876 354680 10928 354686
rect 10876 354622 10928 354628
rect 11704 289876 11756 289882
rect 11704 289818 11756 289824
rect 10876 274712 10928 274718
rect 10876 274654 10928 274660
rect 10784 108996 10836 109002
rect 10784 108938 10836 108944
rect 10600 98864 10652 98870
rect 10600 98806 10652 98812
rect 10506 40080 10562 40089
rect 10506 40015 10562 40024
rect 9496 39704 9548 39710
rect 9496 39646 9548 39652
rect 9404 39228 9456 39234
rect 9404 39170 9456 39176
rect 10888 39166 10916 274654
rect 11716 244254 11744 289818
rect 11704 244248 11756 244254
rect 11704 244190 11756 244196
rect 11704 193248 11756 193254
rect 11704 193190 11756 193196
rect 10966 44568 11022 44577
rect 10966 44503 11022 44512
rect 10876 39160 10928 39166
rect 10876 39102 10928 39108
rect 8944 34400 8996 34406
rect 8944 34342 8996 34348
rect 6656 6886 6868 6914
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 2792 5001 2820 5238
rect 2778 4992 2834 5001
rect 2778 4927 2834 4936
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 20 3188 72 3194
rect 20 3130 72 3136
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 32 480 60 3130
rect 3344 480 3372 3606
rect 6656 480 6684 6886
rect 10980 3534 11008 44503
rect 11716 15162 11744 193190
rect 13096 176662 13124 447102
rect 14476 284306 14504 560254
rect 16500 306338 16528 702406
rect 19720 699718 19748 703520
rect 23032 702434 23060 703520
rect 23032 702406 23428 702434
rect 19708 699712 19760 699718
rect 19708 699654 19760 699660
rect 20628 699712 20680 699718
rect 20628 699654 20680 699660
rect 19984 656940 20036 656946
rect 19984 656882 20036 656888
rect 19996 651438 20024 656882
rect 17960 651432 18012 651438
rect 17960 651374 18012 651380
rect 19984 651432 20036 651438
rect 19984 651374 20036 651380
rect 17972 650026 18000 651374
rect 17880 649998 18000 650026
rect 17880 645930 17908 649998
rect 17868 645924 17920 645930
rect 17868 645866 17920 645872
rect 20260 637356 20312 637362
rect 20260 637298 20312 637304
rect 20272 632126 20300 637298
rect 17224 632120 17276 632126
rect 17224 632062 17276 632068
rect 20260 632120 20312 632126
rect 20260 632062 20312 632068
rect 17236 619614 17264 632062
rect 19156 632052 19208 632058
rect 19156 631994 19208 632000
rect 19168 629678 19196 631994
rect 19156 629672 19208 629678
rect 19156 629614 19208 629620
rect 17960 623892 18012 623898
rect 17960 623834 18012 623840
rect 17972 621058 18000 623834
rect 19984 623824 20036 623830
rect 19984 623766 20036 623772
rect 17880 621030 18000 621058
rect 17224 619608 17276 619614
rect 17224 619550 17276 619556
rect 17880 619546 17908 621030
rect 17868 619540 17920 619546
rect 17868 619482 17920 619488
rect 18052 614168 18104 614174
rect 18052 614110 18104 614116
rect 18064 611182 18092 614110
rect 18788 614100 18840 614106
rect 18788 614042 18840 614048
rect 18052 611176 18104 611182
rect 18052 611118 18104 611124
rect 18800 610026 18828 614042
rect 18788 610020 18840 610026
rect 18788 609962 18840 609968
rect 19996 607170 20024 623766
rect 20076 621036 20128 621042
rect 20076 620978 20128 620984
rect 20088 614174 20116 620978
rect 20076 614168 20128 614174
rect 20076 614110 20128 614116
rect 17960 607164 18012 607170
rect 17960 607106 18012 607112
rect 19984 607164 20036 607170
rect 19984 607106 20036 607112
rect 17972 604654 18000 607106
rect 20168 606756 20220 606762
rect 20168 606698 20220 606704
rect 20180 605130 20208 606698
rect 20168 605124 20220 605130
rect 20168 605066 20220 605072
rect 17960 604648 18012 604654
rect 17960 604590 18012 604596
rect 16488 306332 16540 306338
rect 16488 306274 16540 306280
rect 14464 284300 14516 284306
rect 14464 284242 14516 284248
rect 13084 176656 13136 176662
rect 13084 176598 13136 176604
rect 12072 173868 12124 173874
rect 12072 173810 12124 173816
rect 12084 166598 12112 173810
rect 12072 166592 12124 166598
rect 12072 166534 12124 166540
rect 14464 166592 14516 166598
rect 14464 166534 14516 166540
rect 14476 155922 14504 166534
rect 17868 161492 17920 161498
rect 17868 161434 17920 161440
rect 14464 155916 14516 155922
rect 14464 155858 14516 155864
rect 15200 155916 15252 155922
rect 15200 155858 15252 155864
rect 15212 152114 15240 155858
rect 15200 152108 15252 152114
rect 15200 152050 15252 152056
rect 17224 152108 17276 152114
rect 17224 152050 17276 152056
rect 17236 144906 17264 152050
rect 11796 144900 11848 144906
rect 11796 144842 11848 144848
rect 17224 144900 17276 144906
rect 17224 144842 17276 144848
rect 11808 137562 11836 144842
rect 11796 137556 11848 137562
rect 11796 137498 11848 137504
rect 14464 137556 14516 137562
rect 14464 137498 14516 137504
rect 14476 126954 14504 137498
rect 13084 126948 13136 126954
rect 13084 126890 13136 126896
rect 14464 126948 14516 126954
rect 14464 126890 14516 126896
rect 15200 126948 15252 126954
rect 15200 126890 15252 126896
rect 13096 122262 13124 126890
rect 15212 123214 15240 126890
rect 15844 126880 15896 126886
rect 15844 126822 15896 126828
rect 15200 123208 15252 123214
rect 15200 123150 15252 123156
rect 13084 122256 13136 122262
rect 13084 122198 13136 122204
rect 14372 122256 14424 122262
rect 14372 122198 14424 122204
rect 12440 117360 12492 117366
rect 12440 117302 12492 117308
rect 12452 115802 12480 117302
rect 14384 117298 14412 122198
rect 14372 117292 14424 117298
rect 14372 117234 14424 117240
rect 12440 115796 12492 115802
rect 12440 115738 12492 115744
rect 12440 110424 12492 110430
rect 12440 110366 12492 110372
rect 12452 107642 12480 110366
rect 12440 107636 12492 107642
rect 12440 107578 12492 107584
rect 15856 100026 15884 126822
rect 17224 123208 17276 123214
rect 17224 123150 17276 123156
rect 16212 115796 16264 115802
rect 16212 115738 16264 115744
rect 16224 108322 16252 115738
rect 16212 108316 16264 108322
rect 16212 108258 16264 108264
rect 17236 107574 17264 123150
rect 17316 117292 17368 117298
rect 17316 117234 17368 117240
rect 17328 110498 17356 117234
rect 17316 110492 17368 110498
rect 17316 110434 17368 110440
rect 17408 107636 17460 107642
rect 17408 107578 17460 107584
rect 17224 107568 17276 107574
rect 17224 107510 17276 107516
rect 17420 104854 17448 107578
rect 17408 104848 17460 104854
rect 17408 104790 17460 104796
rect 15844 100020 15896 100026
rect 15844 99962 15896 99968
rect 11796 98864 11848 98870
rect 11796 98806 11848 98812
rect 11808 91934 11836 98806
rect 16488 96620 16540 96626
rect 16488 96562 16540 96568
rect 16500 95146 16528 96562
rect 16500 95118 16620 95146
rect 16592 92546 16620 95118
rect 16580 92540 16632 92546
rect 16580 92482 16632 92488
rect 11796 91928 11848 91934
rect 11796 91870 11848 91876
rect 13728 91928 13780 91934
rect 13728 91870 13780 91876
rect 13740 88398 13768 91870
rect 13728 88392 13780 88398
rect 13728 88334 13780 88340
rect 15200 88324 15252 88330
rect 15200 88266 15252 88272
rect 15212 85610 15240 88266
rect 15200 85604 15252 85610
rect 15200 85546 15252 85552
rect 13728 39364 13780 39370
rect 13728 39306 13780 39312
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 13740 3534 13768 39306
rect 17880 3534 17908 161434
rect 18052 144900 18104 144906
rect 18052 144842 18104 144848
rect 18064 141166 18092 144842
rect 18052 141160 18104 141166
rect 18052 141102 18104 141108
rect 20640 114510 20668 699654
rect 22100 645856 22152 645862
rect 22100 645798 22152 645804
rect 22112 641730 22140 645798
rect 22020 641702 22140 641730
rect 22020 637362 22048 641702
rect 22744 640348 22796 640354
rect 22744 640290 22796 640296
rect 22008 637356 22060 637362
rect 22008 637298 22060 637304
rect 21364 630624 21416 630630
rect 21364 630566 21416 630572
rect 21376 621042 21404 630566
rect 22100 627428 22152 627434
rect 22100 627370 22152 627376
rect 22112 623830 22140 627370
rect 22756 623898 22784 640290
rect 22744 623892 22796 623898
rect 22744 623834 22796 623840
rect 22100 623824 22152 623830
rect 22100 623766 22152 623772
rect 21364 621036 21416 621042
rect 21364 620978 21416 620984
rect 21364 619608 21416 619614
rect 21364 619550 21416 619556
rect 21376 614174 21404 619550
rect 21364 614168 21416 614174
rect 21364 614110 21416 614116
rect 22100 614168 22152 614174
rect 22100 614110 22152 614116
rect 22112 610042 22140 614110
rect 22020 610014 22140 610042
rect 22020 606762 22048 610014
rect 22008 606756 22060 606762
rect 22008 606698 22060 606704
rect 21364 604512 21416 604518
rect 21364 604454 21416 604460
rect 21376 525774 21404 604454
rect 21732 559836 21784 559842
rect 21732 559778 21784 559784
rect 21744 556170 21772 559778
rect 21732 556164 21784 556170
rect 21732 556106 21784 556112
rect 21364 525768 21416 525774
rect 21364 525710 21416 525716
rect 21364 520328 21416 520334
rect 21364 520270 21416 520276
rect 21376 234598 21404 520270
rect 21456 426488 21508 426494
rect 21456 426430 21508 426436
rect 21468 295322 21496 426430
rect 21456 295316 21508 295322
rect 21456 295258 21508 295264
rect 21364 234592 21416 234598
rect 21364 234534 21416 234540
rect 21180 141160 21232 141166
rect 21180 141102 21232 141108
rect 21192 139466 21220 141102
rect 21180 139460 21232 139466
rect 21180 139402 21232 139408
rect 20628 114504 20680 114510
rect 20628 114446 20680 114452
rect 20168 110424 20220 110430
rect 20168 110366 20220 110372
rect 19984 108316 20036 108322
rect 19984 108258 20036 108264
rect 18328 104848 18380 104854
rect 18328 104790 18380 104796
rect 18340 101046 18368 104790
rect 18328 101040 18380 101046
rect 18328 100982 18380 100988
rect 19996 100774 20024 108258
rect 20180 107642 20208 110366
rect 20168 107636 20220 107642
rect 20168 107578 20220 107584
rect 22836 107636 22888 107642
rect 22836 107578 22888 107584
rect 20076 107568 20128 107574
rect 20076 107510 20128 107516
rect 20088 102542 20116 107510
rect 20076 102536 20128 102542
rect 20076 102478 20128 102484
rect 21548 102536 21600 102542
rect 21548 102478 21600 102484
rect 21364 101040 21416 101046
rect 21364 100982 21416 100988
rect 19984 100768 20036 100774
rect 19984 100710 20036 100716
rect 20720 100020 20772 100026
rect 20720 99962 20772 99968
rect 20732 95198 20760 99962
rect 20720 95192 20772 95198
rect 20720 95134 20772 95140
rect 18604 85536 18656 85542
rect 18604 85478 18656 85484
rect 18616 77246 18644 85478
rect 21376 77314 21404 100982
rect 21456 100768 21508 100774
rect 21456 100710 21508 100716
rect 21468 84250 21496 100710
rect 21560 100638 21588 102478
rect 21548 100632 21600 100638
rect 21548 100574 21600 100580
rect 22744 100632 22796 100638
rect 22744 100574 22796 100580
rect 22756 91118 22784 100574
rect 22848 99142 22876 107578
rect 22836 99136 22888 99142
rect 22836 99078 22888 99084
rect 22836 95192 22888 95198
rect 22836 95134 22888 95140
rect 22744 91112 22796 91118
rect 22744 91054 22796 91060
rect 22848 86970 22876 95134
rect 22836 86964 22888 86970
rect 22836 86906 22888 86912
rect 21456 84244 21508 84250
rect 21456 84186 21508 84192
rect 21364 77308 21416 77314
rect 21364 77250 21416 77256
rect 18604 77240 18656 77246
rect 18604 77182 18656 77188
rect 20628 77240 20680 77246
rect 20628 77182 20680 77188
rect 20640 71482 20668 77182
rect 20640 71454 20760 71482
rect 20732 68338 20760 71454
rect 20720 68332 20772 68338
rect 20720 68274 20772 68280
rect 20628 43512 20680 43518
rect 20628 43454 20680 43460
rect 20640 3534 20668 43454
rect 23400 39681 23428 702406
rect 26344 700126 26372 703520
rect 26332 700120 26384 700126
rect 26332 700062 26384 700068
rect 27528 700120 27580 700126
rect 27528 700062 27580 700068
rect 27540 664766 27568 700062
rect 29656 698970 29684 703520
rect 32968 702434 32996 703520
rect 32968 702406 33088 702434
rect 29644 698964 29696 698970
rect 29644 698906 29696 698912
rect 27528 664760 27580 664766
rect 27528 664702 27580 664708
rect 23480 659932 23532 659938
rect 23480 659874 23532 659880
rect 23492 656946 23520 659874
rect 32220 658232 32272 658238
rect 32220 658174 32272 658180
rect 31024 657212 31076 657218
rect 31024 657154 31076 657160
rect 23480 656940 23532 656946
rect 23480 656882 23532 656888
rect 29828 655512 29880 655518
rect 29828 655454 29880 655460
rect 29000 651432 29052 651438
rect 29000 651374 29052 651380
rect 26700 650072 26752 650078
rect 26700 650014 26752 650020
rect 24952 645992 25004 645998
rect 24952 645934 25004 645940
rect 24964 640354 24992 645934
rect 26712 645930 26740 650014
rect 29012 648786 29040 651374
rect 29840 650078 29868 655454
rect 31036 651438 31064 657154
rect 32232 655586 32260 658174
rect 32220 655580 32272 655586
rect 32220 655522 32272 655528
rect 32956 654220 33008 654226
rect 32956 654162 33008 654168
rect 31024 651432 31076 651438
rect 31024 651374 31076 651380
rect 29828 650072 29880 650078
rect 29828 650014 29880 650020
rect 27068 648780 27120 648786
rect 27068 648722 27120 648728
rect 29000 648780 29052 648786
rect 29000 648722 29052 648728
rect 27080 645998 27108 648722
rect 28264 647556 28316 647562
rect 28264 647498 28316 647504
rect 27068 645992 27120 645998
rect 27068 645934 27120 645940
rect 26700 645924 26752 645930
rect 26700 645866 26752 645872
rect 27620 640416 27672 640422
rect 27620 640358 27672 640364
rect 24952 640348 25004 640354
rect 24952 640290 25004 640296
rect 27632 639010 27660 640358
rect 28172 640348 28224 640354
rect 28172 640290 28224 640296
rect 27540 638982 27660 639010
rect 26240 637356 26292 637362
rect 26240 637298 26292 637304
rect 23480 634772 23532 634778
rect 23480 634714 23532 634720
rect 23492 632126 23520 634714
rect 23480 632120 23532 632126
rect 26252 632074 26280 637298
rect 27540 634846 27568 638982
rect 28184 637362 28212 640290
rect 28172 637356 28224 637362
rect 28172 637298 28224 637304
rect 27528 634840 27580 634846
rect 27528 634782 27580 634788
rect 23480 632062 23532 632068
rect 26160 632046 26280 632074
rect 24860 631372 24912 631378
rect 24860 631314 24912 631320
rect 24872 629354 24900 631314
rect 26160 630698 26188 632046
rect 26148 630692 26200 630698
rect 26148 630634 26200 630640
rect 26884 630692 26936 630698
rect 26884 630634 26936 630640
rect 24780 629326 24900 629354
rect 24780 627434 24808 629326
rect 24768 627428 24820 627434
rect 24768 627370 24820 627376
rect 26896 619614 26924 630634
rect 26884 619608 26936 619614
rect 26884 619550 26936 619556
rect 25504 618316 25556 618322
rect 25504 618258 25556 618264
rect 24124 556232 24176 556238
rect 24124 556174 24176 556180
rect 24136 103494 24164 556174
rect 25516 147626 25544 618258
rect 28276 614174 28304 647498
rect 32968 647290 32996 654162
rect 31484 647284 31536 647290
rect 31484 647226 31536 647232
rect 32956 647284 33008 647290
rect 32956 647226 33008 647232
rect 31496 645250 31524 647226
rect 29920 645244 29972 645250
rect 29920 645186 29972 645192
rect 31484 645244 31536 645250
rect 31484 645186 31536 645192
rect 29932 640354 29960 645186
rect 30380 643136 30432 643142
rect 30380 643078 30432 643084
rect 30392 640422 30420 643078
rect 30380 640416 30432 640422
rect 30380 640358 30432 640364
rect 29920 640348 29972 640354
rect 29920 640290 29972 640296
rect 32956 638988 33008 638994
rect 32956 638930 33008 638936
rect 32968 635186 32996 638930
rect 30380 635180 30432 635186
rect 30380 635122 30432 635128
rect 32956 635180 33008 635186
rect 32956 635122 33008 635128
rect 30104 633412 30156 633418
rect 30104 633354 30156 633360
rect 30116 630698 30144 633354
rect 30392 632074 30420 635122
rect 30300 632046 30420 632074
rect 30300 631378 30328 632046
rect 30288 631372 30340 631378
rect 30288 631314 30340 631320
rect 30104 630692 30156 630698
rect 30104 630634 30156 630640
rect 32404 625252 32456 625258
rect 32404 625194 32456 625200
rect 32416 615466 32444 625194
rect 32404 615460 32456 615466
rect 32404 615402 32456 615408
rect 28264 614168 28316 614174
rect 28264 614110 28316 614116
rect 29644 614168 29696 614174
rect 29644 614110 29696 614116
rect 28264 587988 28316 587994
rect 28264 587930 28316 587936
rect 28276 575550 28304 587930
rect 26884 575544 26936 575550
rect 26884 575486 26936 575492
rect 28264 575544 28316 575550
rect 28264 575486 28316 575492
rect 26896 568614 26924 575486
rect 25596 568608 25648 568614
rect 25596 568550 25648 568556
rect 26884 568608 26936 568614
rect 26884 568550 26936 568556
rect 25608 559842 25636 568550
rect 25596 559836 25648 559842
rect 25596 559778 25648 559784
rect 26884 494080 26936 494086
rect 26884 494022 26936 494028
rect 26896 315994 26924 494022
rect 29656 404326 29684 614110
rect 29736 603152 29788 603158
rect 29736 603094 29788 603100
rect 29748 587994 29776 603094
rect 29736 587988 29788 587994
rect 29736 587930 29788 587936
rect 29644 404320 29696 404326
rect 29644 404262 29696 404268
rect 26884 315988 26936 315994
rect 26884 315930 26936 315936
rect 25504 147620 25556 147626
rect 25504 147562 25556 147568
rect 24216 139392 24268 139398
rect 24216 139334 24268 139340
rect 24228 131170 24256 139334
rect 24216 131164 24268 131170
rect 24216 131106 24268 131112
rect 25504 131164 25556 131170
rect 25504 131106 25556 131112
rect 25516 115190 25544 131106
rect 25504 115184 25556 115190
rect 25504 115126 25556 115132
rect 27620 115184 27672 115190
rect 27620 115126 27672 115132
rect 27632 110498 27660 115126
rect 27620 110492 27672 110498
rect 27620 110434 27672 110440
rect 29644 110492 29696 110498
rect 29644 110434 29696 110440
rect 24124 103488 24176 103494
rect 24124 103430 24176 103436
rect 24124 99136 24176 99142
rect 24124 99078 24176 99084
rect 24136 88330 24164 99078
rect 25688 92472 25740 92478
rect 25688 92414 25740 92420
rect 25504 91044 25556 91050
rect 25504 90986 25556 90992
rect 24124 88324 24176 88330
rect 24124 88266 24176 88272
rect 24124 86964 24176 86970
rect 24124 86906 24176 86912
rect 23940 84176 23992 84182
rect 23940 84118 23992 84124
rect 23952 79422 23980 84118
rect 23940 79416 23992 79422
rect 23940 79358 23992 79364
rect 24136 74594 24164 86906
rect 24860 82816 24912 82822
rect 24860 82758 24912 82764
rect 24872 78674 24900 82758
rect 24860 78668 24912 78674
rect 24860 78610 24912 78616
rect 25412 77240 25464 77246
rect 25412 77182 25464 77188
rect 24124 74588 24176 74594
rect 24124 74530 24176 74536
rect 25424 69086 25452 77182
rect 25516 77110 25544 90986
rect 25596 88324 25648 88330
rect 25596 88266 25648 88272
rect 25504 77104 25556 77110
rect 25504 77046 25556 77052
rect 25608 75954 25636 88266
rect 25700 83162 25728 92414
rect 29656 88330 29684 110434
rect 29644 88324 29696 88330
rect 29644 88266 29696 88272
rect 32404 88324 32456 88330
rect 32404 88266 32456 88272
rect 25688 83156 25740 83162
rect 25688 83098 25740 83104
rect 27528 83156 27580 83162
rect 27528 83098 27580 83104
rect 25780 79416 25832 79422
rect 25780 79358 25832 79364
rect 25596 75948 25648 75954
rect 25596 75890 25648 75896
rect 25792 73166 25820 79358
rect 27540 79082 27568 83098
rect 27528 79076 27580 79082
rect 27528 79018 27580 79024
rect 29000 79076 29052 79082
rect 29000 79018 29052 79024
rect 27252 78668 27304 78674
rect 27252 78610 27304 78616
rect 26976 77104 27028 77110
rect 26976 77046 27028 77052
rect 26884 75948 26936 75954
rect 26884 75890 26936 75896
rect 25780 73160 25832 73166
rect 25780 73102 25832 73108
rect 25412 69080 25464 69086
rect 25412 69022 25464 69028
rect 26896 60246 26924 75890
rect 26988 63782 27016 77046
rect 27264 75886 27292 78610
rect 29012 77314 29040 79018
rect 32416 78674 32444 88266
rect 32404 78668 32456 78674
rect 32404 78610 32456 78616
rect 29000 77308 29052 77314
rect 29000 77250 29052 77256
rect 27252 75880 27304 75886
rect 27252 75822 27304 75828
rect 30288 75880 30340 75886
rect 30288 75822 30340 75828
rect 30300 74534 30328 75822
rect 27528 74520 27580 74526
rect 30300 74506 30420 74534
rect 27528 74462 27580 74468
rect 27252 73160 27304 73166
rect 27252 73102 27304 73108
rect 27264 70514 27292 73102
rect 27540 71806 27568 74462
rect 27528 71800 27580 71806
rect 27528 71742 27580 71748
rect 29092 71732 29144 71738
rect 29092 71674 29144 71680
rect 27252 70508 27304 70514
rect 27252 70450 27304 70456
rect 29104 69086 29132 71674
rect 30392 69902 30420 74506
rect 31024 70508 31076 70514
rect 31024 70450 31076 70456
rect 30380 69896 30432 69902
rect 30380 69838 30432 69844
rect 29092 69080 29144 69086
rect 29092 69022 29144 69028
rect 27620 69012 27672 69018
rect 27620 68954 27672 68960
rect 27632 67590 27660 68954
rect 29644 68332 29696 68338
rect 29644 68274 29696 68280
rect 27620 67584 27672 67590
rect 27620 67526 27672 67532
rect 26976 63776 27028 63782
rect 26976 63718 27028 63724
rect 26884 60240 26936 60246
rect 26884 60182 26936 60188
rect 29656 51678 29684 68274
rect 30288 67584 30340 67590
rect 30288 67526 30340 67532
rect 30300 62694 30328 67526
rect 31036 64190 31064 70450
rect 32496 69012 32548 69018
rect 32496 68954 32548 68960
rect 31024 64184 31076 64190
rect 31024 64126 31076 64132
rect 32404 64184 32456 64190
rect 32404 64126 32456 64132
rect 31484 63776 31536 63782
rect 31484 63718 31536 63724
rect 30288 62688 30340 62694
rect 30288 62630 30340 62636
rect 31496 59362 31524 63718
rect 32312 62688 32364 62694
rect 32312 62630 32364 62636
rect 31668 60240 31720 60246
rect 31668 60182 31720 60188
rect 31484 59356 31536 59362
rect 31484 59298 31536 59304
rect 31680 59242 31708 60182
rect 31680 59214 31800 59242
rect 31772 56642 31800 59214
rect 32324 57934 32352 62630
rect 32312 57928 32364 57934
rect 32312 57870 32364 57876
rect 31760 56636 31812 56642
rect 31760 56578 31812 56584
rect 29644 51672 29696 51678
rect 29644 51614 29696 51620
rect 32416 46918 32444 64126
rect 32508 52358 32536 68954
rect 32496 52352 32548 52358
rect 32496 52294 32548 52300
rect 32404 46912 32456 46918
rect 32404 46854 32456 46860
rect 33060 41206 33088 702406
rect 36464 699854 36492 703520
rect 39776 702434 39804 703520
rect 39592 702406 39804 702434
rect 38660 701004 38712 701010
rect 38660 700946 38712 700952
rect 38016 700868 38068 700874
rect 38016 700810 38068 700816
rect 37096 700800 37148 700806
rect 37096 700742 37148 700748
rect 36452 699848 36504 699854
rect 36452 699790 36504 699796
rect 35900 661224 35952 661230
rect 35900 661166 35952 661172
rect 35162 660784 35218 660793
rect 35162 660719 35218 660728
rect 34520 658232 34572 658238
rect 34520 658174 34572 658180
rect 34532 654634 34560 658174
rect 33140 654628 33192 654634
rect 33140 654570 33192 654576
rect 34520 654628 34572 654634
rect 34520 654570 34572 654576
rect 33152 647562 33180 654570
rect 33140 647556 33192 647562
rect 33140 647498 33192 647504
rect 34520 645924 34572 645930
rect 34520 645866 34572 645872
rect 34532 643142 34560 645866
rect 34520 643136 34572 643142
rect 34520 643078 34572 643084
rect 34612 643136 34664 643142
rect 34612 643078 34664 643084
rect 34624 638994 34652 643078
rect 34612 638988 34664 638994
rect 34612 638930 34664 638936
rect 35176 633486 35204 660719
rect 35912 660498 35940 661166
rect 35820 660470 35940 660498
rect 35820 657218 35848 660470
rect 37004 660408 37056 660414
rect 37004 660350 37056 660356
rect 37016 658306 37044 660350
rect 37004 658300 37056 658306
rect 37004 658242 37056 658248
rect 35808 657212 35860 657218
rect 35808 657154 35860 657160
rect 36912 657076 36964 657082
rect 36912 657018 36964 657024
rect 36924 654226 36952 657018
rect 36912 654220 36964 654226
rect 36912 654162 36964 654168
rect 36912 648576 36964 648582
rect 36912 648518 36964 648524
rect 36924 645930 36952 648518
rect 36912 645924 36964 645930
rect 36912 645866 36964 645872
rect 35256 636200 35308 636206
rect 35256 636142 35308 636148
rect 35164 633480 35216 633486
rect 35164 633422 35216 633428
rect 35268 626550 35296 636142
rect 33784 626544 33836 626550
rect 33784 626486 33836 626492
rect 35256 626544 35308 626550
rect 35256 626486 35308 626492
rect 33796 603158 33824 626486
rect 33784 603152 33836 603158
rect 33784 603094 33836 603100
rect 33784 592068 33836 592074
rect 33784 592010 33836 592016
rect 33796 212498 33824 592010
rect 35164 541000 35216 541006
rect 35164 540942 35216 540948
rect 33876 368552 33928 368558
rect 33876 368494 33928 368500
rect 33784 212492 33836 212498
rect 33784 212434 33836 212440
rect 33888 132462 33916 368494
rect 35176 293962 35204 540942
rect 37108 324290 37136 700742
rect 37464 700528 37516 700534
rect 37464 700470 37516 700476
rect 37188 699848 37240 699854
rect 37188 699790 37240 699796
rect 37096 324284 37148 324290
rect 37096 324226 37148 324232
rect 35164 293956 35216 293962
rect 35164 293898 35216 293904
rect 33876 132456 33928 132462
rect 33876 132398 33928 132404
rect 36544 78668 36596 78674
rect 36544 78610 36596 78616
rect 33784 77240 33836 77246
rect 33784 77182 33836 77188
rect 33796 60654 33824 77182
rect 35164 69896 35216 69902
rect 35164 69838 35216 69844
rect 35176 63578 35204 69838
rect 35164 63572 35216 63578
rect 35164 63514 35216 63520
rect 33784 60648 33836 60654
rect 33784 60590 33836 60596
rect 34520 60648 34572 60654
rect 34520 60590 34572 60596
rect 33140 59356 33192 59362
rect 33140 59298 33192 59304
rect 33152 56166 33180 59298
rect 34428 57928 34480 57934
rect 34428 57870 34480 57876
rect 33140 56160 33192 56166
rect 33140 56102 33192 56108
rect 34440 52578 34468 57870
rect 34532 55758 34560 60590
rect 35624 56568 35676 56574
rect 35624 56510 35676 56516
rect 34520 55752 34572 55758
rect 34520 55694 34572 55700
rect 35636 53106 35664 56510
rect 35624 53100 35676 53106
rect 35624 53042 35676 53048
rect 34440 52550 34560 52578
rect 34428 51672 34480 51678
rect 34428 51614 34480 51620
rect 34440 49586 34468 51614
rect 34532 49774 34560 52550
rect 34520 49768 34572 49774
rect 34520 49710 34572 49716
rect 34440 49558 34560 49586
rect 34532 47666 34560 49558
rect 34520 47660 34572 47666
rect 34520 47602 34572 47608
rect 36268 47660 36320 47666
rect 36268 47602 36320 47608
rect 34520 46912 34572 46918
rect 34520 46854 34572 46860
rect 34428 44328 34480 44334
rect 34428 44270 34480 44276
rect 33048 41200 33100 41206
rect 33048 41142 33100 41148
rect 23386 39672 23442 39681
rect 23386 39607 23442 39616
rect 26516 4956 26568 4962
rect 26516 4898 26568 4904
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 9968 480 9996 3470
rect 13280 480 13308 3470
rect 16592 480 16620 3470
rect 19904 480 19932 3470
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23216 480 23244 2994
rect 26528 480 26556 4898
rect 34440 3534 34468 44270
rect 34532 44130 34560 46854
rect 36280 45014 36308 47602
rect 36268 45008 36320 45014
rect 36268 44950 36320 44956
rect 34520 44124 34572 44130
rect 34520 44066 34572 44072
rect 36556 44062 36584 78610
rect 36636 56160 36688 56166
rect 36636 56102 36688 56108
rect 36648 46918 36676 56102
rect 36820 55752 36872 55758
rect 36820 55694 36872 55700
rect 36728 52352 36780 52358
rect 36728 52294 36780 52300
rect 36636 46912 36688 46918
rect 36636 46854 36688 46860
rect 36544 44056 36596 44062
rect 36544 43998 36596 44004
rect 36740 43722 36768 52294
rect 36832 51406 36860 55694
rect 36820 51400 36872 51406
rect 36820 51342 36872 51348
rect 37096 44668 37148 44674
rect 37096 44610 37148 44616
rect 36728 43716 36780 43722
rect 36728 43658 36780 43664
rect 37108 3534 37136 44610
rect 37200 40050 37228 699790
rect 37372 661292 37424 661298
rect 37372 661234 37424 661240
rect 37280 660272 37332 660278
rect 37280 660214 37332 660220
rect 37292 657082 37320 660214
rect 37384 658170 37412 661234
rect 37372 658164 37424 658170
rect 37372 658106 37424 658112
rect 37280 657076 37332 657082
rect 37280 657018 37332 657024
rect 37372 652792 37424 652798
rect 37372 652734 37424 652740
rect 37384 648582 37412 652734
rect 37372 648576 37424 648582
rect 37372 648518 37424 648524
rect 37280 648508 37332 648514
rect 37280 648450 37332 648456
rect 37292 643142 37320 648450
rect 37372 643204 37424 643210
rect 37372 643146 37424 643152
rect 37280 643136 37332 643142
rect 37280 643078 37332 643084
rect 37384 625258 37412 643146
rect 37372 625252 37424 625258
rect 37372 625194 37424 625200
rect 37476 449274 37504 700470
rect 37832 661904 37884 661910
rect 37832 661846 37884 661852
rect 37556 661700 37608 661706
rect 37556 661642 37608 661648
rect 37464 449268 37516 449274
rect 37464 449210 37516 449216
rect 37464 318844 37516 318850
rect 37464 318786 37516 318792
rect 37280 46912 37332 46918
rect 37280 46854 37332 46860
rect 37292 43586 37320 46854
rect 37280 43580 37332 43586
rect 37280 43522 37332 43528
rect 37188 40044 37240 40050
rect 37188 39986 37240 39992
rect 37476 4826 37504 318786
rect 37568 280158 37596 661642
rect 37648 660884 37700 660890
rect 37648 660826 37700 660832
rect 37556 280152 37608 280158
rect 37556 280094 37608 280100
rect 37556 251252 37608 251258
rect 37556 251194 37608 251200
rect 37568 44606 37596 251194
rect 37660 248130 37688 660826
rect 37740 660068 37792 660074
rect 37740 660010 37792 660016
rect 37752 658306 37780 660010
rect 37740 658300 37792 658306
rect 37740 658242 37792 658248
rect 37740 658164 37792 658170
rect 37740 658106 37792 658112
rect 37648 248124 37700 248130
rect 37648 248066 37700 248072
rect 37752 240106 37780 658106
rect 37740 240100 37792 240106
rect 37740 240042 37792 240048
rect 37844 190126 37872 661846
rect 37924 660952 37976 660958
rect 37924 660894 37976 660900
rect 37936 636274 37964 660894
rect 37924 636268 37976 636274
rect 37924 636210 37976 636216
rect 38028 543425 38056 700810
rect 38108 700664 38160 700670
rect 38108 700606 38160 700612
rect 38014 543416 38070 543425
rect 38014 543351 38070 543360
rect 38014 520976 38070 520985
rect 38014 520911 38070 520920
rect 37922 480720 37978 480729
rect 37922 480655 37978 480664
rect 37832 190120 37884 190126
rect 37832 190062 37884 190068
rect 37556 44600 37608 44606
rect 37556 44542 37608 44548
rect 37936 5234 37964 480655
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 38028 3806 38056 520911
rect 38120 122641 38148 700606
rect 38292 700324 38344 700330
rect 38292 700266 38344 700272
rect 38200 660748 38252 660754
rect 38200 660690 38252 660696
rect 38106 122632 38162 122641
rect 38106 122567 38162 122576
rect 38212 68785 38240 660690
rect 38198 68776 38254 68785
rect 38198 68711 38254 68720
rect 38108 63504 38160 63510
rect 38108 63446 38160 63452
rect 38120 52494 38148 63446
rect 38108 52488 38160 52494
rect 38108 52430 38160 52436
rect 38108 51400 38160 51406
rect 38108 51342 38160 51348
rect 38120 44441 38148 51342
rect 38200 49700 38252 49706
rect 38200 49642 38252 49648
rect 38212 44470 38240 49642
rect 38200 44464 38252 44470
rect 38106 44432 38162 44441
rect 38200 44406 38252 44412
rect 38106 44367 38162 44376
rect 38304 38894 38332 700266
rect 38384 699916 38436 699922
rect 38384 699858 38436 699864
rect 38396 39030 38424 699858
rect 38568 665032 38620 665038
rect 38568 664974 38620 664980
rect 38476 663808 38528 663814
rect 38476 663750 38528 663756
rect 38384 39024 38436 39030
rect 38384 38966 38436 38972
rect 38292 38888 38344 38894
rect 38292 38830 38344 38836
rect 38016 3800 38068 3806
rect 38016 3742 38068 3748
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 29828 2916 29880 2922
rect 29828 2858 29880 2864
rect 29840 480 29868 2858
rect 33152 480 33180 3470
rect 36648 480 36676 3470
rect 38488 3330 38516 663750
rect 38580 3942 38608 664974
rect 38672 565729 38700 700946
rect 38844 700596 38896 700602
rect 38844 700538 38896 700544
rect 38752 661020 38804 661026
rect 38752 660962 38804 660968
rect 38764 659841 38792 660962
rect 38750 659832 38806 659841
rect 38750 659767 38806 659776
rect 38856 658442 38884 700538
rect 39488 700256 39540 700262
rect 39488 700198 39540 700204
rect 39212 699984 39264 699990
rect 39212 699926 39264 699932
rect 38936 662312 38988 662318
rect 38936 662254 38988 662260
rect 38844 658436 38896 658442
rect 38844 658378 38896 658384
rect 38948 658186 38976 662254
rect 39028 660476 39080 660482
rect 39028 660418 39080 660424
rect 38764 658158 38976 658186
rect 38658 565720 38714 565729
rect 38658 565655 38714 565664
rect 38660 561672 38712 561678
rect 38660 561614 38712 561620
rect 38672 561377 38700 561614
rect 38658 561368 38714 561377
rect 38658 561303 38714 561312
rect 38658 556880 38714 556889
rect 38658 556815 38714 556824
rect 38672 556238 38700 556815
rect 38660 556232 38712 556238
rect 38660 556174 38712 556180
rect 38660 539572 38712 539578
rect 38660 539514 38712 539520
rect 38672 539073 38700 539514
rect 38658 539064 38714 539073
rect 38658 538999 38714 539008
rect 38660 529984 38712 529990
rect 38658 529952 38660 529961
rect 38712 529952 38714 529961
rect 38658 529887 38714 529896
rect 38660 525768 38712 525774
rect 38660 525710 38712 525716
rect 38672 525473 38700 525710
rect 38658 525464 38714 525473
rect 38658 525399 38714 525408
rect 38658 512136 38714 512145
rect 38658 512071 38714 512080
rect 38568 3936 38620 3942
rect 38568 3878 38620 3884
rect 38476 3324 38528 3330
rect 38476 3266 38528 3272
rect 38672 2854 38700 512071
rect 38764 503169 38792 658158
rect 38844 658096 38896 658102
rect 38844 658038 38896 658044
rect 38856 655489 38884 658038
rect 38936 657212 38988 657218
rect 38936 657154 38988 657160
rect 38842 655480 38898 655489
rect 38842 655415 38898 655424
rect 38844 655376 38896 655382
rect 38844 655318 38896 655324
rect 38856 652798 38884 655318
rect 38844 652792 38896 652798
rect 38844 652734 38896 652740
rect 38844 651364 38896 651370
rect 38844 651306 38896 651312
rect 38856 650865 38884 651306
rect 38842 650856 38898 650865
rect 38842 650791 38898 650800
rect 38844 650752 38896 650758
rect 38844 650694 38896 650700
rect 38856 648514 38884 650694
rect 38844 648508 38896 648514
rect 38844 648450 38896 648456
rect 38844 647216 38896 647222
rect 38844 647158 38896 647164
rect 38856 646513 38884 647158
rect 38842 646504 38898 646513
rect 38842 646439 38898 646448
rect 38948 644474 38976 657154
rect 38856 644446 38976 644474
rect 38856 643210 38884 644446
rect 38844 643204 38896 643210
rect 38844 643146 38896 643152
rect 38844 643068 38896 643074
rect 38844 643010 38896 643016
rect 38856 641889 38884 643010
rect 38842 641880 38898 641889
rect 38842 641815 38898 641824
rect 38934 628416 38990 628425
rect 38934 628351 38990 628360
rect 38842 619440 38898 619449
rect 38842 619375 38898 619384
rect 38856 618322 38884 619375
rect 38844 618316 38896 618322
rect 38844 618258 38896 618264
rect 38842 615088 38898 615097
rect 38842 615023 38898 615032
rect 38856 614174 38884 615023
rect 38844 614168 38896 614174
rect 38844 614110 38896 614116
rect 38844 601656 38896 601662
rect 38842 601624 38844 601633
rect 38896 601624 38898 601633
rect 38842 601559 38898 601568
rect 38844 597508 38896 597514
rect 38844 597450 38896 597456
rect 38856 597281 38884 597450
rect 38842 597272 38898 597281
rect 38842 597207 38898 597216
rect 38842 592512 38898 592521
rect 38842 592447 38898 592456
rect 38856 592074 38884 592447
rect 38844 592068 38896 592074
rect 38844 592010 38896 592016
rect 38844 589280 38896 589286
rect 38844 589222 38896 589228
rect 38856 588305 38884 589222
rect 38842 588296 38898 588305
rect 38842 588231 38898 588240
rect 38948 582894 38976 628351
rect 38936 582888 38988 582894
rect 38936 582830 38988 582836
rect 39040 579329 39068 660418
rect 39120 660136 39172 660142
rect 39120 660078 39172 660084
rect 39026 579320 39082 579329
rect 39026 579255 39082 579264
rect 38842 574560 38898 574569
rect 38842 574495 38898 574504
rect 38856 574122 38884 574495
rect 38844 574116 38896 574122
rect 38844 574058 38896 574064
rect 39132 570353 39160 660078
rect 39118 570344 39174 570353
rect 39118 570279 39174 570288
rect 39120 569016 39172 569022
rect 39120 568958 39172 568964
rect 38750 503160 38806 503169
rect 38750 503095 38806 503104
rect 38752 499520 38804 499526
rect 38752 499462 38804 499468
rect 38764 498817 38792 499462
rect 38750 498808 38806 498817
rect 38750 498743 38806 498752
rect 38750 494184 38806 494193
rect 38750 494119 38806 494128
rect 38764 494086 38792 494119
rect 38752 494080 38804 494086
rect 38752 494022 38804 494028
rect 38750 489696 38806 489705
rect 38750 489631 38806 489640
rect 38764 488578 38792 489631
rect 38752 488572 38804 488578
rect 38752 488514 38804 488520
rect 38752 485784 38804 485790
rect 38752 485726 38804 485732
rect 38764 485217 38792 485726
rect 38750 485208 38806 485217
rect 38750 485143 38806 485152
rect 39132 471889 39160 568958
rect 39224 548049 39252 699926
rect 39304 663400 39356 663406
rect 39304 663342 39356 663348
rect 39316 660822 39344 663342
rect 39304 660816 39356 660822
rect 39304 660758 39356 660764
rect 39394 660648 39450 660657
rect 39304 660612 39356 660618
rect 39394 660583 39450 660592
rect 39304 660554 39356 660560
rect 39316 657393 39344 660554
rect 39302 657384 39358 657393
rect 39302 657319 39358 657328
rect 39304 657280 39356 657286
rect 39304 657222 39356 657228
rect 39210 548040 39266 548049
rect 39210 547975 39266 547984
rect 39118 471880 39174 471889
rect 39118 471815 39174 471824
rect 39316 467265 39344 657222
rect 39302 467256 39358 467265
rect 39302 467191 39358 467200
rect 38752 463684 38804 463690
rect 38752 463626 38804 463632
rect 38764 462913 38792 463626
rect 38750 462904 38806 462913
rect 38750 462839 38806 462848
rect 38752 459536 38804 459542
rect 38752 459478 38804 459484
rect 38764 458289 38792 459478
rect 38750 458280 38806 458289
rect 38750 458215 38806 458224
rect 39304 449268 39356 449274
rect 39304 449210 39356 449216
rect 38750 444816 38806 444825
rect 38750 444751 38806 444760
rect 38764 444446 38792 444751
rect 38752 444440 38804 444446
rect 38752 444382 38804 444388
rect 39316 435985 39344 449210
rect 39302 435976 39358 435985
rect 39302 435911 39358 435920
rect 38752 431928 38804 431934
rect 38752 431870 38804 431876
rect 38764 431633 38792 431870
rect 38750 431624 38806 431633
rect 38750 431559 38806 431568
rect 38750 426864 38806 426873
rect 38750 426799 38806 426808
rect 38764 426494 38792 426799
rect 38752 426488 38804 426494
rect 38752 426430 38804 426436
rect 39408 422657 39436 660583
rect 39500 453937 39528 700198
rect 39592 665922 39620 702406
rect 40040 700936 40092 700942
rect 40040 700878 40092 700884
rect 39948 700460 40000 700466
rect 39948 700402 40000 700408
rect 39672 700392 39724 700398
rect 39672 700334 39724 700340
rect 39580 665916 39632 665922
rect 39580 665858 39632 665864
rect 39580 660204 39632 660210
rect 39580 660146 39632 660152
rect 39486 453928 39542 453937
rect 39486 453863 39542 453872
rect 39488 440292 39540 440298
rect 39488 440234 39540 440240
rect 39394 422648 39450 422657
rect 39394 422583 39450 422592
rect 38750 413536 38806 413545
rect 38750 413471 38806 413480
rect 38764 412690 38792 413471
rect 38752 412684 38804 412690
rect 38752 412626 38804 412632
rect 39396 405952 39448 405958
rect 39396 405894 39448 405900
rect 38750 399936 38806 399945
rect 38750 399871 38806 399880
rect 38764 398886 38792 399871
rect 38752 398880 38804 398886
rect 38752 398822 38804 398828
rect 39408 377777 39436 405894
rect 39394 377768 39450 377777
rect 39394 377703 39450 377712
rect 39394 373280 39450 373289
rect 39394 373215 39450 373224
rect 38750 350704 38806 350713
rect 38750 350639 38806 350648
rect 38764 350606 38792 350639
rect 38752 350600 38804 350606
rect 38752 350542 38804 350548
rect 38750 346488 38806 346497
rect 38750 346423 38752 346432
rect 38804 346423 38806 346432
rect 38752 346394 38804 346400
rect 38750 332752 38806 332761
rect 38750 332687 38806 332696
rect 38764 332654 38792 332687
rect 38752 332648 38804 332654
rect 38752 332590 38804 332596
rect 38752 324284 38804 324290
rect 38752 324226 38804 324232
rect 38764 324193 38792 324226
rect 38750 324184 38806 324193
rect 38750 324119 38806 324128
rect 39302 319424 39358 319433
rect 39302 319359 39358 319368
rect 39316 318850 39344 319359
rect 39304 318844 39356 318850
rect 39304 318786 39356 318792
rect 38750 315072 38806 315081
rect 38750 315007 38806 315016
rect 38764 314702 38792 315007
rect 38752 314696 38804 314702
rect 38752 314638 38804 314644
rect 38750 310584 38806 310593
rect 38750 310519 38752 310528
rect 38804 310519 38806 310528
rect 38752 310490 38804 310496
rect 38752 306332 38804 306338
rect 38752 306274 38804 306280
rect 38764 306241 38792 306274
rect 38750 306232 38806 306241
rect 38750 306167 38806 306176
rect 38752 293956 38804 293962
rect 38752 293898 38804 293904
rect 38764 292641 38792 293898
rect 38750 292632 38806 292641
rect 38750 292567 38806 292576
rect 38752 284300 38804 284306
rect 38752 284242 38804 284248
rect 38764 283665 38792 284242
rect 38750 283656 38806 283665
rect 38750 283591 38806 283600
rect 39304 280152 39356 280158
rect 39304 280094 39356 280100
rect 39316 279313 39344 280094
rect 39302 279304 39358 279313
rect 39302 279239 39358 279248
rect 39408 275398 39436 373215
rect 39396 275392 39448 275398
rect 39396 275334 39448 275340
rect 38752 270496 38804 270502
rect 38752 270438 38804 270444
rect 38764 270337 38792 270438
rect 38750 270328 38806 270337
rect 38750 270263 38806 270272
rect 38750 252240 38806 252249
rect 38750 252175 38806 252184
rect 38764 251258 38792 252175
rect 38752 251252 38804 251258
rect 38752 251194 38804 251200
rect 38844 248124 38896 248130
rect 38844 248066 38896 248072
rect 38856 248033 38884 248066
rect 38842 248024 38898 248033
rect 38842 247959 38898 247968
rect 38752 244248 38804 244254
rect 38752 244190 38804 244196
rect 38764 243409 38792 244190
rect 38750 243400 38806 243409
rect 38750 243335 38806 243344
rect 38752 240100 38804 240106
rect 38752 240042 38804 240048
rect 38764 239057 38792 240042
rect 38750 239048 38806 239057
rect 38750 238983 38806 238992
rect 38752 234592 38804 234598
rect 38752 234534 38804 234540
rect 38764 234433 38792 234534
rect 38750 234424 38806 234433
rect 38750 234359 38806 234368
rect 38750 229936 38806 229945
rect 38750 229871 38806 229880
rect 38764 43858 38792 229871
rect 38842 220960 38898 220969
rect 38842 220895 38898 220904
rect 38856 220862 38884 220895
rect 38844 220856 38896 220862
rect 38844 220798 38896 220804
rect 38844 208344 38896 208350
rect 38844 208286 38896 208292
rect 38856 207777 38884 208286
rect 38842 207768 38898 207777
rect 38842 207703 38898 207712
rect 39500 203153 39528 440234
rect 39592 391105 39620 660146
rect 39684 395729 39712 700334
rect 39856 661088 39908 661094
rect 39856 661030 39908 661036
rect 39764 660000 39816 660006
rect 39764 659942 39816 659948
rect 39776 637537 39804 659942
rect 39762 637528 39818 637537
rect 39762 637463 39818 637472
rect 39762 582448 39818 582457
rect 39762 582383 39818 582392
rect 39670 395720 39726 395729
rect 39670 395655 39726 395664
rect 39578 391096 39634 391105
rect 39578 391031 39634 391040
rect 39578 368656 39634 368665
rect 39578 368591 39634 368600
rect 39592 329798 39620 368591
rect 39670 341728 39726 341737
rect 39670 341663 39726 341672
rect 39580 329792 39632 329798
rect 39580 329734 39632 329740
rect 39578 288144 39634 288153
rect 39578 288079 39634 288088
rect 39486 203144 39542 203153
rect 39486 203079 39542 203088
rect 38842 194032 38898 194041
rect 38842 193967 38898 193976
rect 38856 193254 38884 193967
rect 38844 193248 38896 193254
rect 38844 193190 38896 193196
rect 39488 190120 39540 190126
rect 39488 190062 39540 190068
rect 39500 189825 39528 190062
rect 39486 189816 39542 189825
rect 39486 189751 39542 189760
rect 38842 185056 38898 185065
rect 38842 184991 38898 185000
rect 38856 184958 38884 184991
rect 38844 184952 38896 184958
rect 38844 184894 38896 184900
rect 39118 180840 39174 180849
rect 39118 180775 39174 180784
rect 38844 176656 38896 176662
rect 38844 176598 38896 176604
rect 38856 176225 38884 176598
rect 38842 176216 38898 176225
rect 38842 176151 38898 176160
rect 38844 168360 38896 168366
rect 38844 168302 38896 168308
rect 38856 167249 38884 168302
rect 38842 167240 38898 167249
rect 38842 167175 38898 167184
rect 38842 162752 38898 162761
rect 38842 162687 38898 162696
rect 38856 161498 38884 162687
rect 38844 161492 38896 161498
rect 38844 161434 38896 161440
rect 38934 140448 38990 140457
rect 38934 140383 38990 140392
rect 38844 132456 38896 132462
rect 38844 132398 38896 132404
rect 38856 131617 38884 132398
rect 38842 131608 38898 131617
rect 38842 131543 38898 131552
rect 38844 114504 38896 114510
rect 38844 114446 38896 114452
rect 38856 113665 38884 114446
rect 38842 113656 38898 113665
rect 38842 113591 38898 113600
rect 38842 109032 38898 109041
rect 38842 108967 38844 108976
rect 38896 108967 38898 108976
rect 38844 108938 38896 108944
rect 38948 92070 38976 140383
rect 39132 97986 39160 180775
rect 39486 171728 39542 171737
rect 39486 171663 39542 171672
rect 39302 158128 39358 158137
rect 39302 158063 39358 158072
rect 39210 144800 39266 144809
rect 39210 144735 39266 144744
rect 39120 97980 39172 97986
rect 39120 97922 39172 97928
rect 39026 95568 39082 95577
rect 39026 95503 39082 95512
rect 38936 92064 38988 92070
rect 38936 92006 38988 92012
rect 38934 91216 38990 91225
rect 38934 91151 38990 91160
rect 38842 86592 38898 86601
rect 38842 86527 38898 86536
rect 38856 64802 38884 86527
rect 38844 64796 38896 64802
rect 38844 64738 38896 64744
rect 38842 59664 38898 59673
rect 38842 59599 38898 59608
rect 38856 59430 38884 59599
rect 38844 59424 38896 59430
rect 38844 59366 38896 59372
rect 38844 45008 38896 45014
rect 38844 44950 38896 44956
rect 38856 44033 38884 44950
rect 38842 44024 38898 44033
rect 38842 43959 38898 43968
rect 38752 43852 38804 43858
rect 38752 43794 38804 43800
rect 38948 42362 38976 91151
rect 39040 44198 39068 95503
rect 39118 82240 39174 82249
rect 39118 82175 39174 82184
rect 39028 44192 39080 44198
rect 39028 44134 39080 44140
rect 38936 42356 38988 42362
rect 38936 42298 38988 42304
rect 39132 3738 39160 82175
rect 39224 56574 39252 144735
rect 39212 56568 39264 56574
rect 39212 56510 39264 56516
rect 39212 52488 39264 52494
rect 39212 52430 39264 52436
rect 39224 44266 39252 52430
rect 39212 44260 39264 44266
rect 39212 44202 39264 44208
rect 39316 43994 39344 158063
rect 39394 135824 39450 135833
rect 39394 135759 39450 135768
rect 39304 43988 39356 43994
rect 39304 43930 39356 43936
rect 39408 5098 39436 135759
rect 39500 36582 39528 171663
rect 39488 36576 39540 36582
rect 39488 36518 39540 36524
rect 39592 25566 39620 288079
rect 39684 43926 39712 341663
rect 39776 265985 39804 582383
rect 39762 265976 39818 265985
rect 39762 265911 39818 265920
rect 39868 261361 39896 661030
rect 39960 632913 39988 700402
rect 39946 632904 40002 632913
rect 39946 632839 40002 632848
rect 39948 562352 40000 562358
rect 39948 562294 40000 562300
rect 39960 552401 39988 562294
rect 39946 552392 40002 552401
rect 39946 552327 40002 552336
rect 39948 549024 40000 549030
rect 39948 548966 40000 548972
rect 39960 534449 39988 548966
rect 39946 534440 40002 534449
rect 39946 534375 40002 534384
rect 39948 455388 40000 455394
rect 39948 455330 40000 455336
rect 39960 449313 39988 455330
rect 39946 449304 40002 449313
rect 39946 449239 40002 449248
rect 39854 261352 39910 261361
rect 39854 261287 39910 261296
rect 39762 198792 39818 198801
rect 39762 198727 39818 198736
rect 39672 43920 39724 43926
rect 39672 43862 39724 43868
rect 39776 43790 39804 198727
rect 39946 153776 40002 153785
rect 39946 153711 40002 153720
rect 39960 139534 39988 153711
rect 40052 149569 40080 700878
rect 41880 700732 41932 700738
rect 41880 700674 41932 700680
rect 40408 700188 40460 700194
rect 40408 700130 40460 700136
rect 40132 663196 40184 663202
rect 40132 663138 40184 663144
rect 40144 660550 40172 663138
rect 40224 661428 40276 661434
rect 40224 661370 40276 661376
rect 40132 660544 40184 660550
rect 40132 660486 40184 660492
rect 40132 659796 40184 659802
rect 40132 659738 40184 659744
rect 40144 583681 40172 659738
rect 40130 583672 40186 583681
rect 40130 583607 40186 583616
rect 40236 562358 40264 661370
rect 40316 660952 40368 660958
rect 40316 660894 40368 660900
rect 40328 657218 40356 660894
rect 40316 657212 40368 657218
rect 40316 657154 40368 657160
rect 40316 657076 40368 657082
rect 40316 657018 40368 657024
rect 40224 562352 40276 562358
rect 40224 562294 40276 562300
rect 40130 507376 40186 507385
rect 40130 507311 40186 507320
rect 40038 149560 40094 149569
rect 40038 149495 40094 149504
rect 39948 139528 40000 139534
rect 39948 139470 40000 139476
rect 40038 126848 40094 126857
rect 40038 126783 40094 126792
rect 39854 104544 39910 104553
rect 39854 104479 39910 104488
rect 39868 82686 39896 104479
rect 39946 99920 40002 99929
rect 39946 99855 40002 99864
rect 39856 82680 39908 82686
rect 39856 82622 39908 82628
rect 39960 73710 39988 99855
rect 40052 82414 40080 126783
rect 40040 82408 40092 82414
rect 40040 82350 40092 82356
rect 40038 77616 40094 77625
rect 40038 77551 40094 77560
rect 39948 73704 40000 73710
rect 39948 73646 40000 73652
rect 39854 73264 39910 73273
rect 39854 73199 39910 73208
rect 39764 43784 39816 43790
rect 39764 43726 39816 43732
rect 39580 25560 39632 25566
rect 39580 25502 39632 25508
rect 39868 5438 39896 73199
rect 39946 64288 40002 64297
rect 39946 64223 40002 64232
rect 39960 42090 39988 64223
rect 39948 42084 40000 42090
rect 39948 42026 40000 42032
rect 40052 35222 40080 77551
rect 40144 42430 40172 507311
rect 40222 440464 40278 440473
rect 40222 440399 40278 440408
rect 40132 42424 40184 42430
rect 40132 42366 40184 42372
rect 40040 35216 40092 35222
rect 40040 35158 40092 35164
rect 39856 5432 39908 5438
rect 39856 5374 39908 5380
rect 39396 5092 39448 5098
rect 39396 5034 39448 5040
rect 40236 4010 40264 440399
rect 40328 225457 40356 657018
rect 40420 301617 40448 700130
rect 41604 700120 41656 700126
rect 41604 700062 41656 700068
rect 41236 700052 41288 700058
rect 41236 699994 41288 700000
rect 41052 699848 41104 699854
rect 41052 699790 41104 699796
rect 40592 662380 40644 662386
rect 40592 662322 40644 662328
rect 40500 662176 40552 662182
rect 40500 662118 40552 662124
rect 40406 301608 40462 301617
rect 40406 301543 40462 301552
rect 40406 297120 40462 297129
rect 40406 297055 40462 297064
rect 40314 225448 40370 225457
rect 40314 225383 40370 225392
rect 40314 216336 40370 216345
rect 40314 216271 40370 216280
rect 40328 50658 40356 216271
rect 40316 50652 40368 50658
rect 40316 50594 40368 50600
rect 40316 50516 40368 50522
rect 40316 50458 40368 50464
rect 40328 42498 40356 50458
rect 40316 42492 40368 42498
rect 40316 42434 40368 42440
rect 40224 4004 40276 4010
rect 40224 3946 40276 3952
rect 39120 3732 39172 3738
rect 39120 3674 39172 3680
rect 40420 3262 40448 297055
rect 40512 274689 40540 662118
rect 40604 660414 40632 662322
rect 40684 662244 40736 662250
rect 40684 662186 40736 662192
rect 40592 660408 40644 660414
rect 40592 660350 40644 660356
rect 40592 658708 40644 658714
rect 40592 658650 40644 658656
rect 40604 328545 40632 658650
rect 40696 654134 40724 662186
rect 40776 660544 40828 660550
rect 40776 660486 40828 660492
rect 40958 660512 41014 660521
rect 40788 655246 40816 660486
rect 40958 660447 41014 660456
rect 40868 660408 40920 660414
rect 40868 660350 40920 660356
rect 40776 655240 40828 655246
rect 40776 655182 40828 655188
rect 40696 654106 40816 654134
rect 40684 654016 40736 654022
rect 40684 653958 40736 653964
rect 40696 652798 40724 653958
rect 40684 652792 40736 652798
rect 40684 652734 40736 652740
rect 40684 582888 40736 582894
rect 40684 582830 40736 582836
rect 40590 328536 40646 328545
rect 40590 328471 40646 328480
rect 40498 274680 40554 274689
rect 40498 274615 40554 274624
rect 40498 256864 40554 256873
rect 40498 256799 40554 256808
rect 40512 50402 40540 256799
rect 40590 211984 40646 211993
rect 40590 211919 40646 211928
rect 40604 50522 40632 211919
rect 40592 50516 40644 50522
rect 40592 50458 40644 50464
rect 40512 50374 40632 50402
rect 40500 50312 40552 50318
rect 40500 50254 40552 50260
rect 40512 45626 40540 50254
rect 40500 45620 40552 45626
rect 40500 45562 40552 45568
rect 40498 45520 40554 45529
rect 40498 45455 40554 45464
rect 40512 3466 40540 45455
rect 40604 44538 40632 50374
rect 40592 44532 40644 44538
rect 40592 44474 40644 44480
rect 40592 44396 40644 44402
rect 40592 44338 40644 44344
rect 40604 42226 40632 44338
rect 40592 42220 40644 42226
rect 40592 42162 40644 42168
rect 40696 4078 40724 582830
rect 40788 409057 40816 654106
rect 40880 418033 40908 660350
rect 40972 655382 41000 660447
rect 40960 655376 41012 655382
rect 40960 655318 41012 655324
rect 40960 655240 41012 655246
rect 40960 655182 41012 655188
rect 40866 418024 40922 418033
rect 40866 417959 40922 417968
rect 40774 409048 40830 409057
rect 40774 408983 40830 408992
rect 40972 356017 41000 655182
rect 41064 440298 41092 699790
rect 41144 663264 41196 663270
rect 41144 663206 41196 663212
rect 41156 658714 41184 663206
rect 41144 658708 41196 658714
rect 41144 658650 41196 658656
rect 41144 657416 41196 657422
rect 41144 657358 41196 657364
rect 41052 440292 41104 440298
rect 41052 440234 41104 440240
rect 41052 418192 41104 418198
rect 41052 418134 41104 418140
rect 41064 387297 41092 418134
rect 41156 405958 41184 657358
rect 41248 455394 41276 699994
rect 41328 699780 41380 699786
rect 41328 699722 41380 699728
rect 41340 549030 41368 699722
rect 41420 660816 41472 660822
rect 41420 660758 41472 660764
rect 41432 657422 41460 660758
rect 41510 660376 41566 660385
rect 41510 660311 41566 660320
rect 41420 657416 41472 657422
rect 41420 657358 41472 657364
rect 41420 657280 41472 657286
rect 41420 657222 41472 657228
rect 41432 654158 41460 657222
rect 41420 654152 41472 654158
rect 41420 654094 41472 654100
rect 41524 569022 41552 660311
rect 41512 569016 41564 569022
rect 41512 568958 41564 568964
rect 41328 549024 41380 549030
rect 41328 548966 41380 548972
rect 41616 476785 41644 700062
rect 41788 699712 41840 699718
rect 41788 699654 41840 699660
rect 41696 661360 41748 661366
rect 41696 661302 41748 661308
rect 41708 661026 41736 661302
rect 41696 661020 41748 661026
rect 41696 660962 41748 660968
rect 41694 660104 41750 660113
rect 41694 660039 41750 660048
rect 41602 476776 41658 476785
rect 41602 476711 41658 476720
rect 41236 455388 41288 455394
rect 41236 455330 41288 455336
rect 41708 418198 41736 660039
rect 41696 418192 41748 418198
rect 41696 418134 41748 418140
rect 41144 405952 41196 405958
rect 41144 405894 41196 405900
rect 41050 387288 41106 387297
rect 41050 387223 41106 387232
rect 40958 356008 41014 356017
rect 40958 355943 41014 355952
rect 40776 329792 40828 329798
rect 40776 329734 40828 329740
rect 40684 4072 40736 4078
rect 40684 4014 40736 4020
rect 40788 3874 40816 329734
rect 40868 275392 40920 275398
rect 40868 275334 40920 275340
rect 40776 3868 40828 3874
rect 40776 3810 40828 3816
rect 40500 3460 40552 3466
rect 40500 3402 40552 3408
rect 40408 3256 40460 3262
rect 40408 3198 40460 3204
rect 40880 3194 40908 275334
rect 40960 139528 41012 139534
rect 40960 139470 41012 139476
rect 40972 93566 41000 139470
rect 41144 97980 41196 97986
rect 41144 97922 41196 97928
rect 40960 93560 41012 93566
rect 40960 93502 41012 93508
rect 41052 92064 41104 92070
rect 41052 92006 41104 92012
rect 40960 64796 41012 64802
rect 40960 64738 41012 64744
rect 40972 50726 41000 64738
rect 40960 50720 41012 50726
rect 40960 50662 41012 50668
rect 40958 50144 41014 50153
rect 40958 50079 41014 50088
rect 40972 44470 41000 50079
rect 40960 44464 41012 44470
rect 40960 44406 41012 44412
rect 40960 44192 41012 44198
rect 40960 44134 41012 44140
rect 40972 3398 41000 44134
rect 41064 4146 41092 92006
rect 41156 43246 41184 97922
rect 41604 93560 41656 93566
rect 41604 93502 41656 93508
rect 41328 82680 41380 82686
rect 41328 82622 41380 82628
rect 41236 56568 41288 56574
rect 41236 56510 41288 56516
rect 41144 43240 41196 43246
rect 41144 43182 41196 43188
rect 41052 4140 41104 4146
rect 41052 4082 41104 4088
rect 41248 3602 41276 56510
rect 41340 43178 41368 82622
rect 41512 82408 41564 82414
rect 41512 82350 41564 82356
rect 41420 53100 41472 53106
rect 41420 53042 41472 53048
rect 41432 50862 41460 53042
rect 41420 50856 41472 50862
rect 41420 50798 41472 50804
rect 41420 50720 41472 50726
rect 41420 50662 41472 50668
rect 41432 45762 41460 50662
rect 41420 45756 41472 45762
rect 41420 45698 41472 45704
rect 41420 45620 41472 45626
rect 41420 45562 41472 45568
rect 41328 43172 41380 43178
rect 41328 43114 41380 43120
rect 41432 43110 41460 45562
rect 41524 43382 41552 82350
rect 41616 43654 41644 93502
rect 41696 73704 41748 73710
rect 41696 73646 41748 73652
rect 41604 43648 41656 43654
rect 41604 43590 41656 43596
rect 41512 43376 41564 43382
rect 41512 43318 41564 43324
rect 41420 43104 41472 43110
rect 41420 43046 41472 43052
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40960 3392 41012 3398
rect 40960 3334 41012 3340
rect 40868 3188 40920 3194
rect 40868 3130 40920 3136
rect 41708 3126 41736 73646
rect 41800 45830 41828 699654
rect 41788 45824 41840 45830
rect 41788 45766 41840 45772
rect 41892 45642 41920 700674
rect 43088 699922 43116 703520
rect 43076 699916 43128 699922
rect 43076 699858 43128 699864
rect 46400 699718 46428 703520
rect 49712 702434 49740 703520
rect 49712 702406 49924 702434
rect 46388 699712 46440 699718
rect 46388 699654 46440 699660
rect 49792 665168 49844 665174
rect 49792 665110 49844 665116
rect 46572 665032 46624 665038
rect 46572 664974 46624 664980
rect 43628 663808 43680 663814
rect 43628 663750 43680 663756
rect 43640 662932 43668 663750
rect 46584 662932 46612 664974
rect 49804 662932 49832 665110
rect 49896 662658 49924 702406
rect 53024 699718 53052 703520
rect 56336 700738 56364 703520
rect 56324 700732 56376 700738
rect 56324 700674 56376 700680
rect 54484 699984 54536 699990
rect 59648 699961 59676 703520
rect 62960 700738 62988 703520
rect 62948 700732 63000 700738
rect 62948 700674 63000 700680
rect 54484 699926 54536 699932
rect 59634 699952 59690 699961
rect 53012 699712 53064 699718
rect 53012 699654 53064 699660
rect 53656 699712 53708 699718
rect 53656 699654 53708 699660
rect 52736 665848 52788 665854
rect 52736 665790 52788 665796
rect 52748 662932 52776 665790
rect 53668 663066 53696 699654
rect 54496 665174 54524 699926
rect 59634 699887 59690 699896
rect 66272 699825 66300 703520
rect 66258 699816 66314 699825
rect 66258 699751 66314 699760
rect 69584 699718 69612 703520
rect 73080 701010 73108 703520
rect 73068 701004 73120 701010
rect 73068 700946 73120 700952
rect 73160 701004 73212 701010
rect 73160 700946 73212 700952
rect 73172 700890 73200 700946
rect 73080 700862 73200 700890
rect 73080 699961 73108 700862
rect 73066 699952 73122 699961
rect 73066 699887 73122 699896
rect 76392 699786 76420 703520
rect 79704 702434 79732 703520
rect 79704 702406 80008 702434
rect 76380 699780 76432 699786
rect 76380 699722 76432 699728
rect 77208 699780 77260 699786
rect 77208 699722 77260 699728
rect 66904 699712 66956 699718
rect 66904 699654 66956 699660
rect 69572 699712 69624 699718
rect 69572 699654 69624 699660
rect 70308 699712 70360 699718
rect 70308 699654 70360 699660
rect 60004 698964 60056 698970
rect 60004 698906 60056 698912
rect 59728 675844 59780 675850
rect 59728 675786 59780 675792
rect 59740 666602 59768 675786
rect 57796 666596 57848 666602
rect 57796 666538 57848 666544
rect 59728 666596 59780 666602
rect 59728 666538 59780 666544
rect 57808 666505 57836 666538
rect 57794 666496 57850 666505
rect 57794 666431 57850 666440
rect 54484 665168 54536 665174
rect 54484 665110 54536 665116
rect 60016 665038 60044 698906
rect 64144 697604 64196 697610
rect 64144 697546 64196 697552
rect 64156 687478 64184 697546
rect 62764 687472 62816 687478
rect 62764 687414 62816 687420
rect 64144 687472 64196 687478
rect 64144 687414 64196 687420
rect 62776 679046 62804 687414
rect 61292 679040 61344 679046
rect 61292 678982 61344 678988
rect 62764 679040 62816 679046
rect 62764 678982 62816 678988
rect 61304 675850 61332 678982
rect 61292 675844 61344 675850
rect 61292 675786 61344 675792
rect 66916 666534 66944 699654
rect 68560 698964 68612 698970
rect 68560 698906 68612 698912
rect 68572 697610 68600 698906
rect 68560 697604 68612 697610
rect 68560 697546 68612 697552
rect 64880 666528 64932 666534
rect 64880 666470 64932 666476
rect 66904 666528 66956 666534
rect 66904 666470 66956 666476
rect 60004 665032 60056 665038
rect 60004 664974 60056 664980
rect 61660 664964 61712 664970
rect 61660 664906 61712 664912
rect 55586 664048 55642 664057
rect 55586 663983 55642 663992
rect 58806 664048 58862 664057
rect 58806 663983 58862 663992
rect 53656 663060 53708 663066
rect 53656 663002 53708 663008
rect 55600 662932 55628 663983
rect 58820 662932 58848 663983
rect 59268 663332 59320 663338
rect 59268 663274 59320 663280
rect 49884 662652 49936 662658
rect 49884 662594 49936 662600
rect 59280 662017 59308 663274
rect 61672 662932 61700 664906
rect 64892 662932 64920 666470
rect 70320 664970 70348 699654
rect 70952 666324 71004 666330
rect 70952 666266 71004 666272
rect 70308 664964 70360 664970
rect 70308 664906 70360 664912
rect 70964 662932 70992 666266
rect 73802 664320 73858 664329
rect 73802 664255 73858 664264
rect 73816 662932 73844 664255
rect 77220 663134 77248 699722
rect 79980 666126 80008 702406
rect 83016 699786 83044 703520
rect 86328 699786 86356 703520
rect 83004 699780 83056 699786
rect 83004 699722 83056 699728
rect 86316 699780 86368 699786
rect 86316 699722 86368 699728
rect 86868 699780 86920 699786
rect 86868 699722 86920 699728
rect 79968 666120 80020 666126
rect 79968 666062 80020 666068
rect 86040 665984 86092 665990
rect 86040 665926 86092 665932
rect 79876 664896 79928 664902
rect 79876 664838 79928 664844
rect 77208 663128 77260 663134
rect 77208 663070 77260 663076
rect 79888 662932 79916 664838
rect 83004 664828 83056 664834
rect 83004 664770 83056 664776
rect 83016 662932 83044 664770
rect 86052 662932 86080 665926
rect 86880 665718 86908 699722
rect 86868 665712 86920 665718
rect 86868 665654 86920 665660
rect 89640 664902 89668 703520
rect 92952 700505 92980 703520
rect 92938 700496 92994 700505
rect 92938 700431 92994 700440
rect 95252 665990 95280 703582
rect 96080 703474 96108 703582
rect 96222 703520 96334 704960
rect 99534 703520 99646 704960
rect 102846 703520 102958 704960
rect 106158 703520 106270 704960
rect 109654 703520 109766 704960
rect 112966 703520 113078 704960
rect 116278 703520 116390 704960
rect 119590 703520 119702 704960
rect 122902 703520 123014 704960
rect 125612 703582 126100 703610
rect 96264 703474 96292 703520
rect 96080 703446 96292 703474
rect 99576 699718 99604 703520
rect 102888 699786 102916 703520
rect 106200 699854 106228 703520
rect 109696 702434 109724 703520
rect 109696 702406 109816 702434
rect 106188 699848 106240 699854
rect 106188 699790 106240 699796
rect 102876 699780 102928 699786
rect 102876 699722 102928 699728
rect 109684 699780 109736 699786
rect 109684 699722 109736 699728
rect 99564 699712 99616 699718
rect 99564 699654 99616 699660
rect 98184 666528 98236 666534
rect 98184 666470 98236 666476
rect 95240 665984 95292 665990
rect 95240 665926 95292 665932
rect 89628 664896 89680 664902
rect 89628 664838 89680 664844
rect 89076 664692 89128 664698
rect 89076 664634 89128 664640
rect 89088 662932 89116 664634
rect 98196 662932 98224 666470
rect 101036 665100 101088 665106
rect 101036 665042 101088 665048
rect 107200 665100 107252 665106
rect 107200 665042 107252 665048
rect 101048 662932 101076 665042
rect 104164 665032 104216 665038
rect 104164 664974 104216 664980
rect 104176 662932 104204 664974
rect 107212 662932 107240 665042
rect 109696 664698 109724 699722
rect 109788 696250 109816 702406
rect 113008 699854 113036 703520
rect 116320 700641 116348 703520
rect 116306 700632 116362 700641
rect 116306 700567 116362 700576
rect 112996 699848 113048 699854
rect 112996 699790 113048 699796
rect 119632 699718 119660 703520
rect 122944 699718 122972 703520
rect 119620 699712 119672 699718
rect 119620 699654 119672 699660
rect 122104 699712 122156 699718
rect 122104 699654 122156 699660
rect 122932 699712 122984 699718
rect 122932 699654 122984 699660
rect 124128 699712 124180 699718
rect 124128 699654 124180 699660
rect 109776 696244 109828 696250
rect 109776 696186 109828 696192
rect 122116 666194 122144 699654
rect 122104 666188 122156 666194
rect 122104 666130 122156 666136
rect 124140 666058 124168 699654
rect 124128 666052 124180 666058
rect 124128 665994 124180 666000
rect 113272 665168 113324 665174
rect 113272 665110 113324 665116
rect 109684 664692 109736 664698
rect 109684 664634 109736 664640
rect 113284 662932 113312 665110
rect 119344 664828 119396 664834
rect 119344 664770 119396 664776
rect 119356 662932 119384 664770
rect 125324 664692 125376 664698
rect 125324 664634 125376 664640
rect 122472 663468 122524 663474
rect 122472 663410 122524 663416
rect 122484 662932 122512 663410
rect 125336 662932 125364 664634
rect 95082 662794 95188 662810
rect 95082 662788 95200 662794
rect 95082 662782 95148 662788
rect 95148 662730 95200 662736
rect 77208 662720 77260 662726
rect 59910 662688 59966 662697
rect 67850 662658 68232 662674
rect 77050 662668 77208 662674
rect 110420 662720 110472 662726
rect 77050 662662 77260 662668
rect 110354 662668 110420 662674
rect 116768 662720 116820 662726
rect 110354 662662 110472 662668
rect 116426 662668 116768 662674
rect 116426 662662 116820 662668
rect 67850 662652 68244 662658
rect 67850 662646 68192 662652
rect 59910 662623 59912 662632
rect 59964 662623 59966 662632
rect 59912 662594 59964 662600
rect 77050 662646 77248 662662
rect 110354 662646 110460 662662
rect 116426 662646 116808 662662
rect 68192 662594 68244 662600
rect 125612 662386 125640 703582
rect 126072 703474 126100 703582
rect 126214 703520 126326 704960
rect 129526 703520 129638 704960
rect 132838 703520 132950 704960
rect 136150 703520 136262 704960
rect 139462 703520 139574 704960
rect 142774 703520 142886 704960
rect 146270 703520 146382 704960
rect 149582 703520 149694 704960
rect 152894 703520 153006 704960
rect 156206 703520 156318 704960
rect 159518 703520 159630 704960
rect 162830 703520 162942 704960
rect 166142 703520 166254 704960
rect 169454 703520 169566 704960
rect 172766 703520 172878 704960
rect 175292 703582 175964 703610
rect 126256 703474 126284 703520
rect 126072 703446 126284 703474
rect 129004 699848 129056 699854
rect 129004 699790 129056 699796
rect 129016 664698 129044 699790
rect 129568 698970 129596 703520
rect 132880 699922 132908 703520
rect 136192 702434 136220 703520
rect 136192 702406 136588 702434
rect 132868 699916 132920 699922
rect 132868 699858 132920 699864
rect 129556 698964 129608 698970
rect 129556 698906 129608 698912
rect 135904 696244 135956 696250
rect 135904 696186 135956 696192
rect 134432 665984 134484 665990
rect 134432 665926 134484 665932
rect 129004 664692 129056 664698
rect 129004 664634 129056 664640
rect 131396 663876 131448 663882
rect 131396 663818 131448 663824
rect 131408 662932 131436 663818
rect 134444 662932 134472 665926
rect 135916 665038 135944 696186
rect 136560 666262 136588 702406
rect 139504 700058 139532 703520
rect 139492 700052 139544 700058
rect 139492 699994 139544 700000
rect 142816 699854 142844 703520
rect 146312 700126 146340 703520
rect 149624 700534 149652 703520
rect 149612 700528 149664 700534
rect 149612 700470 149664 700476
rect 146300 700120 146352 700126
rect 146300 700062 146352 700068
rect 152936 700058 152964 703520
rect 156248 702434 156276 703520
rect 155972 702406 156276 702434
rect 152924 700052 152976 700058
rect 152924 699994 152976 700000
rect 150348 699916 150400 699922
rect 150348 699858 150400 699864
rect 142804 699848 142856 699854
rect 142804 699790 142856 699796
rect 136548 666256 136600 666262
rect 136548 666198 136600 666204
rect 146484 666188 146536 666194
rect 146484 666130 146536 666136
rect 135904 665032 135956 665038
rect 135904 664974 135956 664980
rect 140412 665032 140464 665038
rect 140412 664974 140464 664980
rect 137468 664692 137520 664698
rect 137468 664634 137520 664640
rect 137480 662932 137508 664634
rect 140424 662932 140452 664974
rect 143540 664624 143592 664630
rect 143540 664566 143592 664572
rect 142160 663808 142212 663814
rect 142160 663750 142212 663756
rect 142172 663338 142200 663750
rect 142160 663332 142212 663338
rect 142160 663274 142212 663280
rect 143552 662932 143580 664566
rect 146496 662932 146524 666130
rect 150360 663794 150388 699858
rect 152464 699848 152516 699854
rect 152464 699790 152516 699796
rect 152476 664630 152504 699790
rect 152464 664624 152516 664630
rect 152464 664566 152516 664572
rect 150176 663766 150388 663794
rect 152556 663808 152608 663814
rect 150176 662946 150204 663766
rect 152556 663750 152608 663756
rect 149730 662918 150204 662946
rect 152568 662932 152596 663750
rect 155972 662386 156000 702406
rect 159560 699990 159588 703520
rect 162872 700233 162900 703520
rect 166184 700534 166212 703520
rect 166172 700528 166224 700534
rect 166172 700470 166224 700476
rect 162858 700224 162914 700233
rect 162858 700159 162914 700168
rect 169496 700126 169524 703520
rect 169484 700120 169536 700126
rect 169484 700062 169536 700068
rect 159548 699984 159600 699990
rect 159548 699926 159600 699932
rect 172808 699718 172836 703520
rect 172796 699712 172848 699718
rect 172796 699654 172848 699660
rect 173808 699712 173860 699718
rect 173808 699654 173860 699660
rect 171876 676388 171928 676394
rect 171876 676330 171928 676336
rect 171888 673538 171916 676330
rect 166264 673532 166316 673538
rect 166264 673474 166316 673480
rect 171876 673532 171928 673538
rect 171876 673474 171928 673480
rect 161848 666460 161900 666466
rect 161848 666402 161900 666408
rect 161860 662932 161888 666402
rect 164792 666188 164844 666194
rect 164792 666130 164844 666136
rect 164804 662932 164832 666130
rect 125600 662380 125652 662386
rect 125600 662322 125652 662328
rect 155960 662380 156012 662386
rect 155960 662322 156012 662328
rect 158548 662250 158654 662266
rect 158536 662244 158654 662250
rect 158588 662238 158654 662244
rect 158536 662186 158588 662192
rect 128372 662114 128478 662130
rect 128360 662108 128478 662114
rect 128412 662102 128478 662108
rect 155802 662114 155908 662130
rect 155802 662108 155920 662114
rect 155802 662102 155868 662108
rect 128360 662050 128412 662056
rect 155868 662050 155920 662056
rect 59266 662008 59322 662017
rect 92386 662008 92442 662017
rect 92138 661966 92386 661994
rect 59266 661943 59322 661952
rect 92386 661943 92442 661952
rect 166276 661881 166304 673474
rect 167920 665780 167972 665786
rect 167920 665722 167972 665728
rect 167932 662932 167960 665722
rect 170772 664624 170824 664630
rect 170772 664566 170824 664572
rect 170784 662932 170812 664566
rect 173716 664556 173768 664562
rect 173716 664498 173768 664504
rect 173728 662932 173756 664498
rect 173820 663882 173848 699654
rect 175292 676394 175320 703582
rect 175936 703474 175964 703582
rect 176078 703520 176190 704960
rect 179390 703520 179502 704960
rect 182886 703520 182998 704960
rect 186198 703520 186310 704960
rect 189510 703520 189622 704960
rect 192822 703520 192934 704960
rect 196134 703520 196246 704960
rect 199446 703520 199558 704960
rect 202758 703520 202870 704960
rect 206070 703520 206182 704960
rect 209382 703520 209494 704960
rect 212694 703520 212806 704960
rect 216006 703520 216118 704960
rect 219502 703520 219614 704960
rect 222814 703520 222926 704960
rect 226126 703520 226238 704960
rect 229438 703520 229550 704960
rect 232750 703520 232862 704960
rect 236062 703520 236174 704960
rect 239374 703520 239486 704960
rect 241532 703582 242572 703610
rect 176120 703474 176148 703520
rect 175936 703446 176148 703474
rect 175924 700120 175976 700126
rect 175924 700062 175976 700068
rect 175280 676388 175332 676394
rect 175280 676330 175332 676336
rect 175936 673454 175964 700062
rect 179432 699718 179460 703520
rect 182928 699786 182956 703520
rect 180064 699780 180116 699786
rect 180064 699722 180116 699728
rect 182916 699780 182968 699786
rect 182916 699722 182968 699728
rect 179420 699712 179472 699718
rect 179420 699654 179472 699660
rect 175936 673426 176056 673454
rect 176028 664562 176056 673426
rect 180076 665038 180104 699722
rect 180708 699712 180760 699718
rect 180708 699654 180760 699660
rect 176936 665032 176988 665038
rect 176936 664974 176988 664980
rect 180064 665032 180116 665038
rect 180064 664974 180116 664980
rect 176016 664556 176068 664562
rect 176016 664498 176068 664504
rect 173808 663876 173860 663882
rect 173808 663818 173860 663824
rect 176948 662932 176976 664974
rect 180720 664494 180748 699654
rect 182916 664624 182968 664630
rect 182916 664566 182968 664572
rect 180708 664488 180760 664494
rect 180708 664430 180760 664436
rect 182928 662932 182956 664566
rect 186240 664562 186268 703520
rect 189552 700194 189580 703520
rect 192864 702434 192892 703520
rect 192864 702406 193168 702434
rect 189540 700188 189592 700194
rect 189540 700130 189592 700136
rect 193140 665650 193168 702406
rect 196176 699718 196204 703520
rect 199488 699718 199516 703520
rect 202800 700126 202828 703520
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 206112 699922 206140 703520
rect 209424 702434 209452 703520
rect 209424 702406 209728 702434
rect 206100 699916 206152 699922
rect 206100 699858 206152 699864
rect 196164 699712 196216 699718
rect 196164 699654 196216 699660
rect 197268 699712 197320 699718
rect 197268 699654 197320 699660
rect 199476 699712 199528 699718
rect 199476 699654 199528 699660
rect 200028 699712 200080 699718
rect 200028 699654 200080 699660
rect 197280 666398 197308 699654
rect 197268 666392 197320 666398
rect 197268 666334 197320 666340
rect 193128 665644 193180 665650
rect 193128 665586 193180 665592
rect 189080 664692 189132 664698
rect 189080 664634 189132 664640
rect 185860 664556 185912 664562
rect 185860 664498 185912 664504
rect 186228 664556 186280 664562
rect 186228 664498 186280 664504
rect 185872 662932 185900 664498
rect 189092 662932 189120 664634
rect 198004 664556 198056 664562
rect 198004 664498 198056 664504
rect 195060 664420 195112 664426
rect 195060 664362 195112 664368
rect 195072 662932 195100 664362
rect 198016 662932 198044 664498
rect 200040 662114 200068 699654
rect 207204 665712 207256 665718
rect 207204 665654 207256 665660
rect 204076 664012 204128 664018
rect 204076 663954 204128 663960
rect 204088 662932 204116 663954
rect 207216 662932 207244 665654
rect 209700 663338 209728 702406
rect 212736 699718 212764 703520
rect 216048 700262 216076 703520
rect 216036 700256 216088 700262
rect 216036 700198 216088 700204
rect 219544 699718 219572 703520
rect 222856 699718 222884 703520
rect 226168 700097 226196 703520
rect 229480 701049 229508 703520
rect 229466 701040 229522 701049
rect 229466 700975 229522 700984
rect 236104 700262 236132 703520
rect 239416 700942 239444 703520
rect 239404 700936 239456 700942
rect 239404 700878 239456 700884
rect 236092 700256 236144 700262
rect 236092 700198 236144 700204
rect 226154 700088 226210 700097
rect 226154 700023 226210 700032
rect 212724 699712 212776 699718
rect 212724 699654 212776 699660
rect 213828 699712 213880 699718
rect 213828 699654 213880 699660
rect 219532 699712 219584 699718
rect 219532 699654 219584 699660
rect 220728 699712 220780 699718
rect 220728 699654 220780 699660
rect 222844 699712 222896 699718
rect 222844 699654 222896 699660
rect 223488 699712 223540 699718
rect 223488 699654 223540 699660
rect 210240 664556 210292 664562
rect 210240 664498 210292 664504
rect 209688 663332 209740 663338
rect 209688 663274 209740 663280
rect 210252 662932 210280 664498
rect 213184 664012 213236 664018
rect 213184 663954 213236 663960
rect 213196 662932 213224 663954
rect 213840 663474 213868 699654
rect 214656 665236 214708 665242
rect 214656 665178 214708 665184
rect 213828 663468 213880 663474
rect 213828 663410 213880 663416
rect 200028 662108 200080 662114
rect 200028 662050 200080 662056
rect 214668 662017 214696 665178
rect 219164 664964 219216 664970
rect 219164 664906 219216 664912
rect 219176 662932 219204 664906
rect 220740 662250 220768 699654
rect 222108 668160 222160 668166
rect 222108 668102 222160 668108
rect 222120 665242 222148 668102
rect 223500 665718 223528 699654
rect 234528 685160 234580 685166
rect 234528 685102 234580 685108
rect 234540 678298 234568 685102
rect 228364 678292 228416 678298
rect 228364 678234 228416 678240
rect 234528 678292 234580 678298
rect 234528 678234 234580 678240
rect 228376 668166 228404 678234
rect 228364 668160 228416 668166
rect 228364 668102 228416 668108
rect 223488 665712 223540 665718
rect 223488 665654 223540 665660
rect 231308 665644 231360 665650
rect 231308 665586 231360 665592
rect 222108 665236 222160 665242
rect 222108 665178 222160 665184
rect 225236 664760 225288 664766
rect 225236 664702 225288 664708
rect 222384 664080 222436 664086
rect 222384 664022 222436 664028
rect 222396 662932 222424 664022
rect 225248 662932 225276 664702
rect 228364 663808 228416 663814
rect 228364 663750 228416 663756
rect 228376 662932 228404 663750
rect 231320 662932 231348 665586
rect 234528 664964 234580 664970
rect 234528 664906 234580 664912
rect 234540 662932 234568 664906
rect 240506 664456 240562 664465
rect 240506 664391 240562 664400
rect 237470 664184 237526 664193
rect 237470 664119 237526 664128
rect 237484 662932 237512 664119
rect 240520 662932 240548 664391
rect 241532 662318 241560 703582
rect 242544 703474 242572 703582
rect 242686 703520 242798 704960
rect 245998 703520 246110 704960
rect 249310 703520 249422 704960
rect 252622 703520 252734 704960
rect 256118 703520 256230 704960
rect 259430 703520 259542 704960
rect 262742 703520 262854 704960
rect 266054 703520 266166 704960
rect 269366 703520 269478 704960
rect 272678 703520 272790 704960
rect 275990 703520 276102 704960
rect 279302 703520 279414 704960
rect 282614 703520 282726 704960
rect 285926 703520 286038 704960
rect 289238 703520 289350 704960
rect 292734 703520 292846 704960
rect 296046 703520 296158 704960
rect 299358 703520 299470 704960
rect 302670 703520 302782 704960
rect 305012 703582 305868 703610
rect 242728 703474 242756 703520
rect 242544 703446 242756 703474
rect 246040 702434 246068 703520
rect 245764 702406 246068 702434
rect 249352 702434 249380 703520
rect 249352 702406 249748 702434
rect 242164 700256 242216 700262
rect 242164 700198 242216 700204
rect 242176 664766 242204 700198
rect 244924 697604 244976 697610
rect 244924 697546 244976 697552
rect 244936 685166 244964 697546
rect 244924 685160 244976 685166
rect 244924 685102 244976 685108
rect 242164 664760 242216 664766
rect 242164 664702 242216 664708
rect 241520 662312 241572 662318
rect 241520 662254 241572 662260
rect 220728 662244 220780 662250
rect 220728 662186 220780 662192
rect 245764 662182 245792 702406
rect 246580 665712 246632 665718
rect 246580 665654 246632 665660
rect 246592 662932 246620 665654
rect 249720 665038 249748 702406
rect 252664 683114 252692 703520
rect 256160 700194 256188 703520
rect 256148 700188 256200 700194
rect 256148 700130 256200 700136
rect 259472 699718 259500 703520
rect 259460 699712 259512 699718
rect 259460 699654 259512 699660
rect 260748 699712 260800 699718
rect 260748 699654 260800 699660
rect 252572 683086 252692 683114
rect 252572 666534 252600 683086
rect 252560 666528 252612 666534
rect 252560 666470 252612 666476
rect 249708 665032 249760 665038
rect 249708 664974 249760 664980
rect 252560 665032 252612 665038
rect 252560 664974 252612 664980
rect 249524 664352 249576 664358
rect 249524 664294 249576 664300
rect 249536 662932 249564 664294
rect 252572 662932 252600 664974
rect 258540 664760 258592 664766
rect 258540 664702 258592 664708
rect 255686 664320 255742 664329
rect 255686 664255 255742 664264
rect 255700 662932 255728 664255
rect 258552 662932 258580 664702
rect 260760 663678 260788 699654
rect 262784 697610 262812 703520
rect 266096 702434 266124 703520
rect 266096 702406 266308 702434
rect 264980 700052 265032 700058
rect 264980 699994 265032 700000
rect 264992 698698 265020 699994
rect 264980 698692 265032 698698
rect 264980 698634 265032 698640
rect 262772 697604 262824 697610
rect 262772 697546 262824 697552
rect 266280 665038 266308 702406
rect 269408 699718 269436 703520
rect 272720 699718 272748 703520
rect 276032 700874 276060 703520
rect 276020 700868 276072 700874
rect 276020 700810 276072 700816
rect 279344 699718 279372 703520
rect 282656 700262 282684 703520
rect 282644 700256 282696 700262
rect 282644 700198 282696 700204
rect 269396 699712 269448 699718
rect 269396 699654 269448 699660
rect 270408 699712 270460 699718
rect 270408 699654 270460 699660
rect 272708 699712 272760 699718
rect 272708 699654 272760 699660
rect 273168 699712 273220 699718
rect 273168 699654 273220 699660
rect 278780 699712 278832 699718
rect 278780 699654 278832 699660
rect 279332 699712 279384 699718
rect 279332 699654 279384 699660
rect 267004 698692 267056 698698
rect 267004 698634 267056 698640
rect 267016 686526 267044 698634
rect 267004 686520 267056 686526
rect 267004 686462 267056 686468
rect 270420 666534 270448 699654
rect 270408 666528 270460 666534
rect 270408 666470 270460 666476
rect 266268 665032 266320 665038
rect 266268 664974 266320 664980
rect 270684 664896 270736 664902
rect 270684 664838 270736 664844
rect 264704 664352 264756 664358
rect 264704 664294 264756 664300
rect 260748 663672 260800 663678
rect 260748 663614 260800 663620
rect 261760 663604 261812 663610
rect 261760 663546 261812 663552
rect 261772 662932 261800 663546
rect 264716 662932 264744 664294
rect 267740 664284 267792 664290
rect 267740 664226 267792 664232
rect 267752 662932 267780 664226
rect 270696 662932 270724 664838
rect 273180 664766 273208 699654
rect 273260 686520 273312 686526
rect 273260 686462 273312 686468
rect 273272 684554 273300 686462
rect 273260 684548 273312 684554
rect 273260 684490 273312 684496
rect 276756 665032 276808 665038
rect 276756 664974 276808 664980
rect 273168 664760 273220 664766
rect 273168 664702 273220 664708
rect 273902 664592 273958 664601
rect 273902 664527 273958 664536
rect 273916 662932 273944 664527
rect 276768 662932 276796 664974
rect 278792 662946 278820 699654
rect 285968 697610 285996 703520
rect 289280 699718 289308 703520
rect 289268 699712 289320 699718
rect 289268 699654 289320 699660
rect 289728 699712 289780 699718
rect 289728 699654 289780 699660
rect 285956 697604 286008 697610
rect 285956 697546 286008 697552
rect 278872 684480 278924 684486
rect 278872 684422 278924 684428
rect 278884 681766 278912 684422
rect 278872 681760 278924 681766
rect 278872 681702 278924 681708
rect 280804 681760 280856 681766
rect 280804 681702 280856 681708
rect 280816 672110 280844 681702
rect 280804 672104 280856 672110
rect 280804 672046 280856 672052
rect 282920 672036 282972 672042
rect 282920 671978 282972 671984
rect 282932 668642 282960 671978
rect 282920 668636 282972 668642
rect 282920 668578 282972 668584
rect 284944 668636 284996 668642
rect 284944 668578 284996 668584
rect 282920 664760 282972 664766
rect 282920 664702 282972 664708
rect 278792 662918 279910 662946
rect 282932 662932 282960 664702
rect 245752 662176 245804 662182
rect 284956 662153 284984 668578
rect 289740 664902 289768 699654
rect 292776 683114 292804 703520
rect 299400 700874 299428 703520
rect 302712 700942 302740 703520
rect 302700 700936 302752 700942
rect 302700 700878 302752 700884
rect 299388 700868 299440 700874
rect 299388 700810 299440 700816
rect 294604 697604 294656 697610
rect 294604 697546 294656 697552
rect 294616 692782 294644 697546
rect 294604 692776 294656 692782
rect 294604 692718 294656 692724
rect 298008 692776 298060 692782
rect 298008 692718 298060 692724
rect 298020 689042 298048 692718
rect 298008 689036 298060 689042
rect 298008 688978 298060 688984
rect 292592 683086 292804 683114
rect 292592 666330 292620 683086
rect 292580 666324 292632 666330
rect 292580 666266 292632 666272
rect 305012 665038 305040 703582
rect 305840 703474 305868 703582
rect 305982 703520 306094 704960
rect 309294 703520 309406 704960
rect 312606 703520 312718 704960
rect 315918 703520 316030 704960
rect 318812 703582 319116 703610
rect 306024 703474 306052 703520
rect 305840 703446 306052 703474
rect 309336 699718 309364 703520
rect 312648 700806 312676 703520
rect 315960 703050 315988 703520
rect 314660 703044 314712 703050
rect 314660 702986 314712 702992
rect 315948 703044 316000 703050
rect 315948 702986 316000 702992
rect 312636 700800 312688 700806
rect 312636 700742 312688 700748
rect 309324 699712 309376 699718
rect 309324 699654 309376 699660
rect 310428 699712 310480 699718
rect 310428 699654 310480 699660
rect 305092 689036 305144 689042
rect 305092 688978 305144 688984
rect 305104 685166 305132 688978
rect 305092 685160 305144 685166
rect 305092 685102 305144 685108
rect 310244 685160 310296 685166
rect 310244 685102 310296 685108
rect 310256 682650 310284 685102
rect 310244 682644 310296 682650
rect 310244 682586 310296 682592
rect 304080 665032 304132 665038
rect 304080 664974 304132 664980
rect 305000 665032 305052 665038
rect 305000 664974 305052 664980
rect 289728 664896 289780 664902
rect 289728 664838 289780 664844
rect 295062 664728 295118 664737
rect 295062 664663 295118 664672
rect 288900 664216 288952 664222
rect 288900 664158 288952 664164
rect 291936 664216 291988 664222
rect 291936 664158 291988 664164
rect 288912 662932 288940 664158
rect 291948 662932 291976 664158
rect 295076 662932 295104 664663
rect 304092 662932 304120 664974
rect 307206 663912 307262 663921
rect 307206 663847 307262 663856
rect 307220 662932 307248 663847
rect 310440 662318 310468 699654
rect 314672 664834 314700 702986
rect 318708 682644 318760 682650
rect 318708 682586 318760 682592
rect 318720 679658 318748 682586
rect 318708 679652 318760 679658
rect 318708 679594 318760 679600
rect 316224 666324 316276 666330
rect 316224 666266 316276 666272
rect 314660 664828 314712 664834
rect 314660 664770 314712 664776
rect 313280 664148 313332 664154
rect 313280 664090 313332 664096
rect 313292 662932 313320 664090
rect 316236 662932 316264 666266
rect 318812 665786 318840 703582
rect 319088 703474 319116 703582
rect 319230 703520 319342 704960
rect 322542 703520 322654 704960
rect 325854 703520 325966 704960
rect 329350 703520 329462 704960
rect 332662 703520 332774 704960
rect 335974 703520 336086 704960
rect 339286 703520 339398 704960
rect 342272 703582 342484 703610
rect 319272 703474 319300 703520
rect 319088 703446 319300 703474
rect 322584 699961 322612 703520
rect 324320 700188 324372 700194
rect 324320 700130 324372 700136
rect 325608 700188 325660 700194
rect 325608 700130 325660 700136
rect 322570 699952 322626 699961
rect 322570 699887 322626 699896
rect 324332 696250 324360 700130
rect 324320 696244 324372 696250
rect 324320 696186 324372 696192
rect 318800 665780 318852 665786
rect 318800 665722 318852 665728
rect 322296 664284 322348 664290
rect 322296 664226 322348 664232
rect 319352 664148 319404 664154
rect 319352 664090 319404 664096
rect 319364 662932 319392 664090
rect 322308 662932 322336 664226
rect 325620 662946 325648 700130
rect 325896 683114 325924 703520
rect 329392 700806 329420 703520
rect 329380 700800 329432 700806
rect 329380 700742 329432 700748
rect 326804 700120 326856 700126
rect 326804 700062 326856 700068
rect 326816 699650 326844 700062
rect 332704 699825 332732 703520
rect 336016 700670 336044 703520
rect 339328 702434 339356 703520
rect 339328 702406 339448 702434
rect 336004 700664 336056 700670
rect 336004 700606 336056 700612
rect 332690 699816 332746 699825
rect 332690 699751 332746 699760
rect 326804 699644 326856 699650
rect 326804 699586 326856 699592
rect 334624 699644 334676 699650
rect 334624 699586 334676 699592
rect 331864 696244 331916 696250
rect 331864 696186 331916 696192
rect 331876 690062 331904 696186
rect 334636 692646 334664 699586
rect 334624 692640 334676 692646
rect 334624 692582 334676 692588
rect 336464 692640 336516 692646
rect 336464 692582 336516 692588
rect 331864 690056 331916 690062
rect 331864 689998 331916 690004
rect 333244 690056 333296 690062
rect 333244 689998 333296 690004
rect 325712 683086 325924 683114
rect 325712 666466 325740 683086
rect 333256 680950 333284 689998
rect 336476 689790 336504 692582
rect 336464 689784 336516 689790
rect 336464 689726 336516 689732
rect 338764 689784 338816 689790
rect 338764 689726 338816 689732
rect 338776 681766 338804 689726
rect 338764 681760 338816 681766
rect 338764 681702 338816 681708
rect 333244 680944 333296 680950
rect 333244 680886 333296 680892
rect 333980 680944 334032 680950
rect 333980 680886 334032 680892
rect 332508 680400 332560 680406
rect 332508 680342 332560 680348
rect 331864 679652 331916 679658
rect 331864 679594 331916 679600
rect 331876 671362 331904 679594
rect 331864 671356 331916 671362
rect 331864 671298 331916 671304
rect 325700 666460 325752 666466
rect 325700 666402 325752 666408
rect 332520 665038 332548 680342
rect 333992 676870 334020 680886
rect 333980 676864 334032 676870
rect 333980 676806 334032 676812
rect 331312 665032 331364 665038
rect 331312 664974 331364 664980
rect 332508 665032 332560 665038
rect 332508 664974 332560 664980
rect 337384 665032 337436 665038
rect 337384 664974 337436 664980
rect 328276 663536 328328 663542
rect 328276 663478 328328 663484
rect 325450 662918 325648 662946
rect 328288 662932 328316 663478
rect 331324 662932 331352 664974
rect 334440 664760 334492 664766
rect 334440 664702 334492 664708
rect 334452 662932 334480 664702
rect 336740 664420 336792 664426
rect 336740 664362 336792 664368
rect 336752 663746 336780 664362
rect 336740 663740 336792 663746
rect 336740 663682 336792 663688
rect 337396 662932 337424 664974
rect 339420 663542 339448 702406
rect 340144 681760 340196 681766
rect 340144 681702 340196 681708
rect 340156 669390 340184 681702
rect 341524 676864 341576 676870
rect 341524 676806 341576 676812
rect 341536 672586 341564 676806
rect 341524 672580 341576 672586
rect 341524 672522 341576 672528
rect 340144 669384 340196 669390
rect 340144 669326 340196 669332
rect 340512 666460 340564 666466
rect 340512 666402 340564 666408
rect 339408 663536 339460 663542
rect 339408 663478 339460 663484
rect 340524 662932 340552 666402
rect 342272 665038 342300 703582
rect 342456 703474 342484 703582
rect 342598 703520 342710 704960
rect 345910 703520 346022 704960
rect 349222 703520 349334 704960
rect 352534 703520 352646 704960
rect 355846 703520 355958 704960
rect 359158 703520 359270 704960
rect 362470 703520 362582 704960
rect 365966 703520 366078 704960
rect 368492 703582 369164 703610
rect 342640 703474 342668 703520
rect 342456 703446 342668 703474
rect 345952 700670 345980 703520
rect 345940 700664 345992 700670
rect 345940 700606 345992 700612
rect 349264 699825 349292 703520
rect 352472 700732 352524 700738
rect 352472 700674 352524 700680
rect 349250 699816 349306 699825
rect 349250 699751 349306 699760
rect 352484 692774 352512 700674
rect 352576 699718 352604 703520
rect 355888 702434 355916 703520
rect 355888 702406 356008 702434
rect 352748 700732 352800 700738
rect 352748 700674 352800 700680
rect 352656 700120 352708 700126
rect 352656 700062 352708 700068
rect 352564 699712 352616 699718
rect 352564 699654 352616 699660
rect 352484 692746 352604 692774
rect 346308 672580 346360 672586
rect 346308 672522 346360 672528
rect 343640 671356 343692 671362
rect 343640 671298 343692 671304
rect 343652 668545 343680 671298
rect 346124 669248 346176 669254
rect 346124 669190 346176 669196
rect 346320 669202 346348 672522
rect 343638 668536 343694 668545
rect 343638 668471 343694 668480
rect 346136 666505 346164 669190
rect 346320 669174 346440 669202
rect 346122 666496 346178 666505
rect 346122 666431 346178 666440
rect 346412 665786 346440 669174
rect 346400 665780 346452 665786
rect 346400 665722 346452 665728
rect 349068 665780 349120 665786
rect 349068 665722 349120 665728
rect 342260 665032 342312 665038
rect 342260 664974 342312 664980
rect 343454 664456 343510 664465
rect 343454 664391 343510 664400
rect 343468 662932 343496 664391
rect 349080 663794 349108 665722
rect 352576 664834 352604 692746
rect 352668 664970 352696 700062
rect 352760 666466 352788 700674
rect 353208 699712 353260 699718
rect 353208 699654 353260 699660
rect 353220 666466 353248 699654
rect 352748 666460 352800 666466
rect 352748 666402 352800 666408
rect 353208 666460 353260 666466
rect 353208 666402 353260 666408
rect 352656 664964 352708 664970
rect 352656 664906 352708 664912
rect 352564 664828 352616 664834
rect 352564 664770 352616 664776
rect 349528 664352 349580 664358
rect 349528 664294 349580 664300
rect 349080 663785 349200 663794
rect 349080 663776 349214 663785
rect 349080 663766 349158 663776
rect 349158 663711 349214 663720
rect 349540 662932 349568 664294
rect 355980 663746 356008 702406
rect 362512 700602 362540 703520
rect 362500 700596 362552 700602
rect 362500 700538 362552 700544
rect 366008 699825 366036 703520
rect 365994 699816 366050 699825
rect 365994 699751 366050 699760
rect 358636 666256 358688 666262
rect 358636 666198 358688 666204
rect 353300 663740 353352 663746
rect 353300 663682 353352 663688
rect 355968 663740 356020 663746
rect 355968 663682 356020 663688
rect 353312 662425 353340 663682
rect 358648 662932 358676 666198
rect 368492 664970 368520 703582
rect 369136 703474 369164 703582
rect 369278 703520 369390 704960
rect 372590 703520 372702 704960
rect 375392 703582 375788 703610
rect 369320 703474 369348 703520
rect 369136 703446 369348 703474
rect 361672 664964 361724 664970
rect 361672 664906 361724 664912
rect 368480 664964 368532 664970
rect 368480 664906 368532 664912
rect 361684 662932 361712 664906
rect 370688 664420 370740 664426
rect 370688 664362 370740 664368
rect 364800 663808 364852 663814
rect 364800 663750 364852 663756
rect 364812 662932 364840 663750
rect 370700 662932 370728 664362
rect 372632 663406 372660 703520
rect 373816 665032 373868 665038
rect 373816 664974 373868 664980
rect 372620 663400 372672 663406
rect 372620 663342 372672 663348
rect 373828 662932 373856 664974
rect 375392 664426 375420 703582
rect 375760 703474 375788 703582
rect 375902 703520 376014 704960
rect 378152 703582 379100 703610
rect 375944 703474 375972 703520
rect 375760 703446 375972 703474
rect 375380 664420 375432 664426
rect 375380 664362 375432 664368
rect 376760 664420 376812 664426
rect 376760 664362 376812 664368
rect 376772 662932 376800 664362
rect 378152 663270 378180 703582
rect 379072 703474 379100 703582
rect 379214 703520 379326 704960
rect 382526 703520 382638 704960
rect 385838 703520 385950 704960
rect 389150 703520 389262 704960
rect 391952 703582 392348 703610
rect 379256 703474 379284 703520
rect 379072 703446 379284 703474
rect 382568 700126 382596 703520
rect 385880 700738 385908 703520
rect 385868 700732 385920 700738
rect 385868 700674 385920 700680
rect 382556 700120 382608 700126
rect 382556 700062 382608 700068
rect 388812 666528 388864 666534
rect 388812 666470 388864 666476
rect 385960 664964 386012 664970
rect 385960 664906 386012 664912
rect 382740 663944 382792 663950
rect 382740 663886 382792 663892
rect 378140 663264 378192 663270
rect 378140 663206 378192 663212
rect 382752 662932 382780 663886
rect 385972 662932 386000 664906
rect 388824 662932 388852 666470
rect 389192 665038 389220 703520
rect 389180 665032 389232 665038
rect 389180 664974 389232 664980
rect 391952 664426 391980 703582
rect 392320 703474 392348 703582
rect 392462 703520 392574 704960
rect 395774 703520 395886 704960
rect 399086 703520 399198 704960
rect 401612 703582 402468 703610
rect 392504 703474 392532 703520
rect 392320 703446 392532 703474
rect 395816 700602 395844 703520
rect 399128 700913 399156 703520
rect 399114 700904 399170 700913
rect 399114 700839 399170 700848
rect 398748 700732 398800 700738
rect 398748 700674 398800 700680
rect 395804 700596 395856 700602
rect 395804 700538 395856 700544
rect 391940 664420 391992 664426
rect 391940 664362 391992 664368
rect 398760 663794 398788 700674
rect 401612 664970 401640 703582
rect 402440 703474 402468 703582
rect 402582 703520 402694 704960
rect 405894 703520 406006 704960
rect 409206 703520 409318 704960
rect 412518 703520 412630 704960
rect 415830 703520 415942 704960
rect 419142 703520 419254 704960
rect 422454 703520 422566 704960
rect 425766 703520 425878 704960
rect 429078 703520 429190 704960
rect 432390 703520 432502 704960
rect 434732 703582 435588 703610
rect 402624 703474 402652 703520
rect 402440 703446 402652 703474
rect 407120 666392 407172 666398
rect 407120 666334 407172 666340
rect 401600 664964 401652 664970
rect 401600 664906 401652 664912
rect 398576 663766 398788 663794
rect 398576 662946 398604 663766
rect 398130 662918 398604 662946
rect 403716 662992 403768 662998
rect 403768 662940 404110 662946
rect 403716 662934 404110 662940
rect 403728 662918 404110 662934
rect 407132 662932 407160 666334
rect 409892 662930 409998 662946
rect 409880 662924 409998 662930
rect 409932 662918 409998 662924
rect 409880 662866 409932 662872
rect 353298 662416 353354 662425
rect 353298 662351 353354 662360
rect 354036 662380 354088 662386
rect 354036 662322 354088 662328
rect 358268 662380 358320 662386
rect 358268 662322 358320 662328
rect 310428 662312 310480 662318
rect 310428 662254 310480 662260
rect 286416 662176 286468 662182
rect 245752 662118 245804 662124
rect 284942 662144 284998 662153
rect 286074 662124 286416 662130
rect 354048 662153 354076 662322
rect 358280 662153 358308 662322
rect 286074 662118 286468 662124
rect 297822 662144 297878 662153
rect 286074 662102 286456 662118
rect 284942 662079 284998 662088
rect 301410 662144 301466 662153
rect 297878 662102 297942 662130
rect 301162 662102 301410 662130
rect 297822 662079 297878 662088
rect 301410 662079 301466 662088
rect 354034 662144 354090 662153
rect 354034 662079 354090 662088
rect 358266 662144 358322 662153
rect 358266 662079 358322 662088
rect 309692 662040 309744 662046
rect 214654 662008 214710 662017
rect 200776 661978 201158 661994
rect 200764 661972 201158 661978
rect 200816 661966 201158 661972
rect 243910 662008 243966 662017
rect 216338 661978 216628 661994
rect 216338 661972 216640 661978
rect 216338 661966 216588 661972
rect 214654 661943 214710 661952
rect 200764 661914 200816 661920
rect 243570 661966 243910 661994
rect 346952 662040 347004 662046
rect 309744 661988 310086 661994
rect 309692 661982 310086 661988
rect 309704 661966 310086 661982
rect 346610 661988 346952 661994
rect 353022 662008 353078 662017
rect 346610 661982 347004 661988
rect 346610 661966 346992 661982
rect 352682 661966 353022 661994
rect 243910 661943 243966 661952
rect 353022 661943 353078 661952
rect 216588 661914 216640 661920
rect 166262 661872 166318 661881
rect 166262 661807 166318 661816
rect 179510 661872 179566 661881
rect 192390 661872 192446 661881
rect 179566 661830 179814 661858
rect 192050 661830 192390 661858
rect 179510 661807 179566 661816
rect 355966 661872 356022 661881
rect 355626 661830 355966 661858
rect 192390 661807 192446 661816
rect 355966 661807 356022 661816
rect 367282 661872 367338 661881
rect 394790 661872 394846 661881
rect 367338 661830 367678 661858
rect 379532 661842 379822 661858
rect 379520 661836 379822 661842
rect 367282 661807 367338 661816
rect 379572 661830 379822 661836
rect 392058 661842 392440 661858
rect 392058 661836 392452 661842
rect 392058 661830 392400 661836
rect 379520 661778 379572 661784
rect 394846 661830 394910 661858
rect 394790 661807 394846 661816
rect 392400 661778 392452 661784
rect 412560 661774 412588 703520
rect 415872 700738 415900 703520
rect 419184 700738 419212 703520
rect 415860 700732 415912 700738
rect 415860 700674 415912 700680
rect 419172 700732 419224 700738
rect 419172 700674 419224 700680
rect 422496 700466 422524 703520
rect 422484 700460 422536 700466
rect 422484 700402 422536 700408
rect 416044 700120 416096 700126
rect 416044 700062 416096 700068
rect 416056 665038 416084 700062
rect 425808 699990 425836 703520
rect 429120 700126 429148 703520
rect 432432 700398 432460 703520
rect 432420 700392 432472 700398
rect 432420 700334 432472 700340
rect 429108 700120 429160 700126
rect 429108 700062 429160 700068
rect 425796 699984 425848 699990
rect 425796 699926 425848 699932
rect 426348 699984 426400 699990
rect 426348 699926 426400 699932
rect 422208 666256 422260 666262
rect 422208 666198 422260 666204
rect 413192 665032 413244 665038
rect 413192 664974 413244 664980
rect 416044 665032 416096 665038
rect 416044 664974 416096 664980
rect 413204 662932 413232 664974
rect 416136 664420 416188 664426
rect 416136 664362 416188 664368
rect 416148 662932 416176 664362
rect 422220 662932 422248 666198
rect 418804 662856 418856 662862
rect 418856 662804 419198 662810
rect 418804 662798 419198 662804
rect 418816 662782 419198 662798
rect 425072 662386 425270 662402
rect 426360 662386 426388 699926
rect 428188 666460 428240 666466
rect 428188 666402 428240 666408
rect 428200 662932 428228 666402
rect 431316 666120 431368 666126
rect 431316 666062 431368 666068
rect 431328 662932 431356 666062
rect 434732 663202 434760 703582
rect 435560 703474 435588 703582
rect 435702 703520 435814 704960
rect 439198 703520 439310 704960
rect 441632 703582 442396 703610
rect 435744 703474 435772 703520
rect 435560 703446 435772 703474
rect 439240 699718 439268 703520
rect 436744 699712 436796 699718
rect 436744 699654 436796 699660
rect 439228 699712 439280 699718
rect 439228 699654 439280 699660
rect 436756 666262 436784 699654
rect 441632 666330 441660 703582
rect 442368 703474 442396 703582
rect 442510 703520 442622 704960
rect 445822 703520 445934 704960
rect 449134 703520 449246 704960
rect 452446 703520 452558 704960
rect 455758 703520 455870 704960
rect 458192 703582 458956 703610
rect 442552 703474 442580 703520
rect 442368 703446 442580 703474
rect 449176 700777 449204 703520
rect 449162 700768 449218 700777
rect 449162 700703 449218 700712
rect 452488 700233 452516 703520
rect 455800 700466 455828 703520
rect 455788 700460 455840 700466
rect 455788 700402 455840 700408
rect 452474 700224 452530 700233
rect 452474 700159 452530 700168
rect 441620 666324 441672 666330
rect 441620 666266 441672 666272
rect 436744 666256 436796 666262
rect 436744 666198 436796 666204
rect 443460 664828 443512 664834
rect 443460 664770 443512 664776
rect 446496 664828 446548 664834
rect 446496 664770 446548 664776
rect 437478 664320 437534 664329
rect 437478 664255 437534 664264
rect 434720 663196 434772 663202
rect 434720 663138 434772 663144
rect 437492 662932 437520 664255
rect 443472 662932 443500 664770
rect 446508 662932 446536 664770
rect 458192 664698 458220 703582
rect 458928 703474 458956 703582
rect 459070 703520 459182 704960
rect 462382 703520 462494 704960
rect 465694 703520 465806 704960
rect 469006 703520 469118 704960
rect 471992 703582 472204 703610
rect 459112 703474 459140 703520
rect 458928 703446 459140 703474
rect 459468 700392 459520 700398
rect 459468 700334 459520 700340
rect 459480 665038 459508 700334
rect 462424 700194 462452 703520
rect 462412 700188 462464 700194
rect 462412 700130 462464 700136
rect 464988 700188 465040 700194
rect 464988 700130 465040 700136
rect 461584 700120 461636 700126
rect 461584 700062 461636 700068
rect 458640 665032 458692 665038
rect 458640 664974 458692 664980
rect 459468 665032 459520 665038
rect 459468 664974 459520 664980
rect 458180 664692 458232 664698
rect 458180 664634 458232 664640
rect 455512 664624 455564 664630
rect 455512 664566 455564 664572
rect 449346 663912 449402 663921
rect 449346 663847 449402 663856
rect 449360 662932 449388 663847
rect 455524 662932 455552 664566
rect 458652 662932 458680 664974
rect 461596 664630 461624 700062
rect 461584 664624 461636 664630
rect 461584 664566 461636 664572
rect 465000 662946 465028 700130
rect 465736 699718 465764 703520
rect 469048 699825 469076 703520
rect 469034 699816 469090 699825
rect 469034 699751 469090 699760
rect 465724 699712 465776 699718
rect 465724 699654 465776 699660
rect 466368 699712 466420 699718
rect 466368 699654 466420 699660
rect 466380 664970 466408 699654
rect 466368 664964 466420 664970
rect 466368 664906 466420 664912
rect 470692 664896 470744 664902
rect 470692 664838 470744 664844
rect 464738 662918 465028 662946
rect 470704 662932 470732 664838
rect 433892 662856 433944 662862
rect 433944 662804 434286 662810
rect 433892 662798 434286 662804
rect 433904 662782 434286 662798
rect 425060 662380 425270 662386
rect 425112 662374 425270 662380
rect 426348 662380 426400 662386
rect 425060 662322 425112 662328
rect 426348 662322 426400 662328
rect 471992 661910 472020 703582
rect 472176 703474 472204 703582
rect 472318 703520 472430 704960
rect 475814 703520 475926 704960
rect 479126 703520 479238 704960
rect 481652 703582 482324 703610
rect 472360 703474 472388 703520
rect 472176 703446 472388 703474
rect 475856 702434 475884 703520
rect 475856 702406 476068 702434
rect 473728 665032 473780 665038
rect 473728 664974 473780 664980
rect 473740 662932 473768 664974
rect 476040 661910 476068 702406
rect 479168 700126 479196 703520
rect 479156 700120 479208 700126
rect 479156 700062 479208 700068
rect 481652 666194 481680 703582
rect 482296 703474 482324 703582
rect 482438 703520 482550 704960
rect 485750 703520 485862 704960
rect 489062 703520 489174 704960
rect 491312 703582 492260 703610
rect 482480 703474 482508 703520
rect 482296 703446 482508 703474
rect 485792 700126 485820 703520
rect 485780 700120 485832 700126
rect 485780 700062 485832 700068
rect 489104 699825 489132 703520
rect 489184 700052 489236 700058
rect 489184 699994 489236 700000
rect 489090 699816 489146 699825
rect 489090 699751 489146 699760
rect 481640 666188 481692 666194
rect 481640 666130 481692 666136
rect 489196 665038 489224 699994
rect 489184 665032 489236 665038
rect 489184 664974 489236 664980
rect 482928 664896 482980 664902
rect 482928 664838 482980 664844
rect 476856 664692 476908 664698
rect 476856 664634 476908 664640
rect 476868 662932 476896 664634
rect 482940 662932 482968 664838
rect 485872 664624 485924 664630
rect 485872 664566 485924 664572
rect 485884 662932 485912 664566
rect 491312 663814 491340 703582
rect 492232 703474 492260 703582
rect 492374 703520 492486 704960
rect 495686 703520 495798 704960
rect 498998 703520 499110 704960
rect 502310 703520 502422 704960
rect 505622 703520 505734 704960
rect 508934 703520 509046 704960
rect 512012 703582 512316 703610
rect 492416 703474 492444 703520
rect 492232 703446 492444 703474
rect 495728 700330 495756 703520
rect 495716 700324 495768 700330
rect 495716 700266 495768 700272
rect 491944 700256 491996 700262
rect 491944 700198 491996 700204
rect 491956 665038 491984 700198
rect 499040 700058 499068 703520
rect 502352 700913 502380 703520
rect 502338 700904 502394 700913
rect 502338 700839 502394 700848
rect 499028 700052 499080 700058
rect 499028 699994 499080 700000
rect 505664 699718 505692 703520
rect 508976 700330 509004 703520
rect 508964 700324 509016 700330
rect 508964 700266 509016 700272
rect 505652 699712 505704 699718
rect 505652 699654 505704 699660
rect 506388 699712 506440 699718
rect 506388 699654 506440 699660
rect 492220 666120 492272 666126
rect 492220 666062 492272 666068
rect 491944 665032 491996 665038
rect 491944 664974 491996 664980
rect 488816 663808 488868 663814
rect 488816 663750 488868 663756
rect 491300 663808 491352 663814
rect 491300 663750 491352 663756
rect 488828 662932 488856 663750
rect 492232 662946 492260 666062
rect 500960 665032 501012 665038
rect 500960 664974 501012 664980
rect 494796 663876 494848 663882
rect 494796 663818 494848 663824
rect 491970 662918 492260 662946
rect 494808 662932 494836 663818
rect 500972 662932 501000 664974
rect 503994 664864 504050 664873
rect 503994 664799 504050 664808
rect 504008 662932 504036 664799
rect 479340 662856 479392 662862
rect 479392 662804 479734 662810
rect 479340 662798 479734 662804
rect 479352 662782 479734 662798
rect 506400 662590 506428 699654
rect 509884 698352 509936 698358
rect 509884 698294 509936 698300
rect 509896 665038 509924 698294
rect 510068 666052 510120 666058
rect 510068 665994 510120 666000
rect 509884 665032 509936 665038
rect 509884 664974 509936 664980
rect 507032 663876 507084 663882
rect 507032 663818 507084 663824
rect 507044 662932 507072 663818
rect 510080 662932 510108 665994
rect 497556 662584 497608 662590
rect 506388 662584 506440 662590
rect 497608 662532 497950 662538
rect 497556 662526 497950 662532
rect 506388 662526 506440 662532
rect 497568 662510 497950 662526
rect 471980 661904 472032 661910
rect 440238 661872 440294 661881
rect 452106 661872 452162 661881
rect 440294 661830 440358 661858
rect 440238 661807 440294 661816
rect 461122 661872 461178 661881
rect 452162 661830 452502 661858
rect 452106 661807 452162 661816
rect 467194 661872 467250 661881
rect 461178 661830 461518 661858
rect 461122 661807 461178 661816
rect 467250 661830 467590 661858
rect 471980 661846 472032 661852
rect 476028 661904 476080 661910
rect 476028 661846 476080 661852
rect 467194 661807 467250 661816
rect 400588 661768 400640 661774
rect 412548 661768 412600 661774
rect 400640 661716 400982 661722
rect 400588 661710 400982 661716
rect 412548 661710 412600 661716
rect 400600 661694 400982 661710
rect 512012 661706 512040 703582
rect 512288 703474 512316 703582
rect 512430 703520 512542 704960
rect 515742 703520 515854 704960
rect 519054 703520 519166 704960
rect 521672 703582 522252 703610
rect 512472 703474 512500 703520
rect 512288 703446 512500 703474
rect 515784 699718 515812 703520
rect 519096 699718 519124 703520
rect 512644 699712 512696 699718
rect 512644 699654 512696 699660
rect 515772 699712 515824 699718
rect 515772 699654 515824 699660
rect 519084 699712 519136 699718
rect 519084 699654 519136 699660
rect 520188 699712 520240 699718
rect 520188 699654 520240 699660
rect 512656 666126 512684 699654
rect 512644 666120 512696 666126
rect 512644 666062 512696 666068
rect 519084 665916 519136 665922
rect 519084 665858 519136 665864
rect 516140 665032 516192 665038
rect 516140 664974 516192 664980
rect 516152 662932 516180 664974
rect 519096 662932 519124 665858
rect 512642 661736 512698 661745
rect 512000 661700 512052 661706
rect 515218 661736 515274 661745
rect 512698 661694 513038 661722
rect 520200 661706 520228 699654
rect 521672 664766 521700 703582
rect 522224 703474 522252 703582
rect 522366 703520 522478 704960
rect 525678 703520 525790 704960
rect 528572 703582 528876 703610
rect 522408 703474 522436 703520
rect 522224 703446 522436 703474
rect 521660 664760 521712 664766
rect 521660 664702 521712 664708
rect 522304 664760 522356 664766
rect 522304 664702 522356 664708
rect 522316 662932 522344 664702
rect 528190 663912 528246 663921
rect 528190 663847 528246 663856
rect 528204 662932 528232 663847
rect 528572 661881 528600 703582
rect 528848 703474 528876 703582
rect 528990 703520 529102 704960
rect 531332 703582 532188 703610
rect 529032 703474 529060 703520
rect 528848 703446 529060 703474
rect 531332 665990 531360 703582
rect 532160 703474 532188 703582
rect 532302 703520 532414 704960
rect 535614 703520 535726 704960
rect 538926 703520 539038 704960
rect 542238 703520 542350 704960
rect 545550 703520 545662 704960
rect 547892 703582 548932 703610
rect 532344 703474 532372 703520
rect 532160 703446 532372 703474
rect 535656 700194 535684 703520
rect 535644 700188 535696 700194
rect 535644 700130 535696 700136
rect 538968 699825 538996 703520
rect 542280 702434 542308 703520
rect 545592 702434 545620 703520
rect 542096 702406 542308 702434
rect 545316 702406 545620 702434
rect 541992 700868 542044 700874
rect 541992 700810 542044 700816
rect 538954 699816 539010 699825
rect 538954 699751 539010 699760
rect 531320 665984 531372 665990
rect 531320 665926 531372 665932
rect 539600 665168 539652 665174
rect 539600 665110 539652 665116
rect 531320 664964 531372 664970
rect 531320 664906 531372 664912
rect 531332 662932 531360 664906
rect 534172 664488 534224 664494
rect 534172 664430 534224 664436
rect 537392 664488 537444 664494
rect 537392 664430 537444 664436
rect 534184 662932 534212 664430
rect 537404 662932 537432 664430
rect 528558 661872 528614 661881
rect 528558 661807 528614 661816
rect 524786 661736 524842 661745
rect 512642 661671 512698 661680
rect 515218 661671 515220 661680
rect 512000 661642 512052 661648
rect 515272 661671 515274 661680
rect 520188 661700 520240 661706
rect 515220 661642 515272 661648
rect 524842 661694 525182 661722
rect 539612 661706 539640 665110
rect 540336 663808 540388 663814
rect 540336 663750 540388 663756
rect 540348 662932 540376 663750
rect 539600 661700 539652 661706
rect 524786 661671 524842 661680
rect 520188 661642 520240 661648
rect 539600 661642 539652 661648
rect 541898 661600 541954 661609
rect 541898 661535 541954 661544
rect 541912 660890 541940 661535
rect 541900 660884 541952 660890
rect 541900 660826 541952 660832
rect 541900 660748 541952 660754
rect 541900 660690 541952 660696
rect 541912 654294 541940 660690
rect 541900 654288 541952 654294
rect 541900 654230 541952 654236
rect 541900 654146 541952 654152
rect 541900 654088 541952 654094
rect 541912 331022 541940 654088
rect 542004 610881 542032 700810
rect 542096 700369 542124 702406
rect 543924 700936 543976 700942
rect 543924 700878 543976 700884
rect 543832 700800 543884 700806
rect 543832 700742 543884 700748
rect 542268 700732 542320 700738
rect 542268 700674 542320 700680
rect 542176 700460 542228 700466
rect 542176 700402 542228 700408
rect 542082 700360 542138 700369
rect 542082 700295 542138 700304
rect 542084 661224 542136 661230
rect 542084 661166 542136 661172
rect 542096 660929 542124 661166
rect 542082 660920 542138 660929
rect 542082 660855 542138 660864
rect 542084 660272 542136 660278
rect 542084 660214 542136 660220
rect 542096 654242 542124 660214
rect 542188 654362 542216 700402
rect 542280 661366 542308 700674
rect 543740 700664 543792 700670
rect 543740 700606 543792 700612
rect 543648 700596 543700 700602
rect 543648 700538 543700 700544
rect 542820 700528 542872 700534
rect 542820 700470 542872 700476
rect 542360 664828 542412 664834
rect 542360 664770 542412 664776
rect 542268 661360 542320 661366
rect 542268 661302 542320 661308
rect 542268 660816 542320 660822
rect 542268 660758 542320 660764
rect 542176 654356 542228 654362
rect 542176 654298 542228 654304
rect 542096 654214 542216 654242
rect 542084 654152 542136 654158
rect 542084 654094 542136 654100
rect 541990 610872 542046 610881
rect 541990 610807 542046 610816
rect 542096 505986 542124 654094
rect 542188 543250 542216 654214
rect 542280 620362 542308 660758
rect 542268 620356 542320 620362
rect 542268 620298 542320 620304
rect 542176 543244 542228 543250
rect 542176 543186 542228 543192
rect 542084 505980 542136 505986
rect 542084 505922 542136 505928
rect 541990 471880 542046 471889
rect 541990 471815 542046 471824
rect 542004 466313 542032 471815
rect 541990 466304 542046 466313
rect 541990 466239 542046 466248
rect 541990 442504 542046 442513
rect 541990 442439 542046 442448
rect 542004 438977 542032 442439
rect 542082 439104 542138 439113
rect 542082 439039 542138 439048
rect 541990 438968 542046 438977
rect 541990 438903 542046 438912
rect 542096 438161 542124 439039
rect 542082 438152 542138 438161
rect 542082 438087 542138 438096
rect 541900 331016 541952 331022
rect 541900 330958 541952 330964
rect 541898 193352 541954 193361
rect 541898 193287 541954 193296
rect 41800 45614 41920 45642
rect 41800 39982 41828 45614
rect 41880 45566 41932 45572
rect 41880 45508 41932 45514
rect 41892 44305 41920 45508
rect 41878 44296 41934 44305
rect 41878 44231 41934 44240
rect 41880 44192 41932 44198
rect 41880 44134 41932 44140
rect 41892 43314 41920 44134
rect 541912 43586 541940 193287
rect 541990 143984 542046 143993
rect 541990 143919 542046 143928
rect 541900 43580 541952 43586
rect 541900 43522 541952 43528
rect 41880 43308 41932 43314
rect 41880 43250 41932 43256
rect 41880 43036 41932 43042
rect 41880 42978 41932 42984
rect 41788 39976 41840 39982
rect 41788 39918 41840 39924
rect 41892 38758 41920 42978
rect 196072 42424 196124 42430
rect 59266 42392 59322 42401
rect 379428 42424 379480 42430
rect 223946 42392 224002 42401
rect 196072 42366 196124 42372
rect 59266 42327 59322 42336
rect 59280 41392 59308 42327
rect 68006 42256 68062 42265
rect 68006 42191 68062 42200
rect 64892 41534 66102 41562
rect 59280 41364 59400 41392
rect 41984 39778 42012 41140
rect 41972 39772 42024 39778
rect 41972 39714 42024 39720
rect 44088 38956 44140 38962
rect 44088 38898 44140 38904
rect 41880 38752 41932 38758
rect 41880 38694 41932 38700
rect 44100 3534 44128 38898
rect 44928 38690 44956 41140
rect 47872 38894 47900 41140
rect 51092 40050 51120 41140
rect 51080 40044 51132 40050
rect 51080 39986 51132 39992
rect 53944 39370 53972 41140
rect 57178 41126 57928 41154
rect 53932 39364 53984 39370
rect 53932 39306 53984 39312
rect 47860 38888 47912 38894
rect 47860 38830 47912 38836
rect 44916 38684 44968 38690
rect 44916 38626 44968 38632
rect 57900 5506 57928 41126
rect 59372 39370 59400 41364
rect 60108 39817 60136 41140
rect 62132 41126 63158 41154
rect 60094 39808 60150 39817
rect 60094 39743 60150 39752
rect 59360 39364 59412 39370
rect 59360 39306 59412 39312
rect 61384 39364 61436 39370
rect 61384 39306 61436 39312
rect 61396 17950 61424 39306
rect 61384 17944 61436 17950
rect 61384 17886 61436 17892
rect 57888 5500 57940 5506
rect 57888 5442 57940 5448
rect 49884 4888 49936 4894
rect 49884 4830 49936 4836
rect 46572 3800 46624 3806
rect 46572 3742 46624 3748
rect 43260 3528 43312 3534
rect 43260 3470 43312 3476
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 41696 3120 41748 3126
rect 41696 3062 41748 3068
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 39960 480 39988 2926
rect 43272 480 43300 3470
rect 46584 480 46612 3742
rect 49896 480 49924 4830
rect 59820 3800 59872 3806
rect 59820 3742 59872 3748
rect 56506 3496 56562 3505
rect 56506 3431 56562 3440
rect 53196 2848 53248 2854
rect 53196 2790 53248 2796
rect 53208 480 53236 2790
rect 56520 480 56548 3431
rect 59832 480 59860 3742
rect 62132 2922 62160 41126
rect 64512 17944 64564 17950
rect 64512 17886 64564 17892
rect 64524 10334 64552 17886
rect 64512 10328 64564 10334
rect 64512 10270 64564 10276
rect 64892 3058 64920 41534
rect 65984 41404 66036 41410
rect 65984 41346 66036 41352
rect 65996 39778 66024 41346
rect 68020 40526 68048 42191
rect 169668 42152 169720 42158
rect 157430 42120 157486 42129
rect 169668 42094 169720 42100
rect 157430 42055 157486 42064
rect 157444 41410 157472 42055
rect 162872 41410 163070 41426
rect 157432 41404 157484 41410
rect 157432 41346 157484 41352
rect 162860 41404 163070 41410
rect 162912 41398 163070 41404
rect 162860 41346 162912 41352
rect 71780 41336 71832 41342
rect 71832 41284 72174 41290
rect 71780 41278 72174 41284
rect 71792 41262 72174 41278
rect 156616 41274 156998 41290
rect 156604 41268 156998 41274
rect 156656 41262 156998 41268
rect 156604 41210 156656 41216
rect 69216 40662 69244 41140
rect 69204 40656 69256 40662
rect 69204 40598 69256 40604
rect 68008 40520 68060 40526
rect 68008 40462 68060 40468
rect 65984 39772 66036 39778
rect 65984 39714 66036 39720
rect 75288 38758 75316 41140
rect 77312 41126 78246 41154
rect 75276 38752 75328 38758
rect 75276 38694 75328 38700
rect 69664 10328 69716 10334
rect 69664 10270 69716 10276
rect 69676 5030 69704 10270
rect 69756 5364 69808 5370
rect 69756 5306 69808 5312
rect 69664 5024 69716 5030
rect 69664 4966 69716 4972
rect 64880 3052 64932 3058
rect 64880 2994 64932 3000
rect 62120 2916 62172 2922
rect 62120 2858 62172 2864
rect 63132 2916 63184 2922
rect 63132 2858 63184 2864
rect 63144 480 63172 2858
rect 69768 480 69796 5306
rect 73250 3632 73306 3641
rect 73250 3567 73306 3576
rect 73264 480 73292 3567
rect 76564 3052 76616 3058
rect 76564 2994 76616 3000
rect 76576 480 76604 2994
rect 77312 2990 77340 41126
rect 81176 38962 81204 41140
rect 84304 39545 84332 41140
rect 86972 41126 87262 41154
rect 84290 39536 84346 39545
rect 84290 39471 84346 39480
rect 86868 39364 86920 39370
rect 86868 39306 86920 39312
rect 81164 38956 81216 38962
rect 81164 38898 81216 38904
rect 86880 6914 86908 39306
rect 86512 6886 86908 6914
rect 83186 6216 83242 6225
rect 83186 6151 83242 6160
rect 79876 5296 79928 5302
rect 79876 5238 79928 5244
rect 77300 2984 77352 2990
rect 77300 2926 77352 2932
rect 79888 480 79916 5238
rect 83200 480 83228 6151
rect 86512 480 86540 6886
rect 86972 2854 87000 41126
rect 90468 38894 90496 41140
rect 92584 41126 93334 41154
rect 90456 38888 90508 38894
rect 90456 38830 90508 38836
rect 89812 2984 89864 2990
rect 89812 2926 89864 2932
rect 86960 2848 87012 2854
rect 86960 2790 87012 2796
rect 89824 480 89852 2926
rect 92584 2922 92612 41126
rect 96448 40458 96476 41140
rect 96436 40452 96488 40458
rect 96436 40394 96488 40400
rect 93124 6180 93176 6186
rect 93124 6122 93176 6128
rect 92572 2916 92624 2922
rect 92572 2858 92624 2864
rect 93136 480 93164 6122
rect 96434 4856 96490 4865
rect 96434 4791 96490 4800
rect 96448 480 96476 4791
rect 99392 3670 99420 41140
rect 102612 40458 102640 41140
rect 102600 40452 102652 40458
rect 102600 40394 102652 40400
rect 105556 38962 105584 41140
rect 105544 38956 105596 38962
rect 105544 38898 105596 38904
rect 108684 38690 108712 41140
rect 111642 41126 111748 41154
rect 108672 38684 108724 38690
rect 108672 38626 108724 38632
rect 99746 5400 99802 5409
rect 99746 5335 99802 5344
rect 99380 3664 99432 3670
rect 99380 3606 99432 3612
rect 99760 480 99788 5335
rect 111720 4758 111748 41126
rect 114664 38826 114692 41140
rect 117608 39370 117636 41140
rect 120092 41126 120566 41154
rect 117596 39364 117648 39370
rect 117596 39306 117648 39312
rect 114652 38820 114704 38826
rect 114652 38762 114704 38768
rect 119988 38820 120040 38826
rect 119988 38762 120040 38768
rect 120000 6914 120028 38762
rect 119816 6886 120028 6914
rect 111708 4752 111760 4758
rect 111708 4694 111760 4700
rect 116490 3768 116546 3777
rect 116490 3703 116546 3712
rect 113180 3664 113232 3670
rect 113180 3606 113232 3612
rect 106370 3496 106426 3505
rect 106370 3431 106426 3440
rect 103060 3120 103112 3126
rect 103060 3062 103112 3068
rect 103072 480 103100 3062
rect 106384 480 106412 3431
rect 113192 480 113220 3606
rect 116504 480 116532 3703
rect 119816 480 119844 6886
rect 120092 2990 120120 41126
rect 123772 40050 123800 41140
rect 123760 40044 123812 40050
rect 123760 39986 123812 39992
rect 126716 39370 126744 41140
rect 126704 39364 126756 39370
rect 126704 39306 126756 39312
rect 129844 38758 129872 41140
rect 132696 39953 132724 41140
rect 135824 40526 135852 41140
rect 138860 40526 138888 41140
rect 140792 41126 141910 41154
rect 135812 40520 135864 40526
rect 135812 40462 135864 40468
rect 138848 40520 138900 40526
rect 138848 40462 138900 40468
rect 132682 39944 132738 39953
rect 132682 39879 132738 39888
rect 131764 38888 131816 38894
rect 131764 38830 131816 38836
rect 131856 38888 131908 38894
rect 131856 38830 131908 38836
rect 129832 38752 129884 38758
rect 129832 38694 129884 38700
rect 131028 38752 131080 38758
rect 131028 38694 131080 38700
rect 126428 5024 126480 5030
rect 126428 4966 126480 4972
rect 129740 5024 129792 5030
rect 129740 4966 129792 4972
rect 120080 2984 120132 2990
rect 120080 2926 120132 2932
rect 123116 2984 123168 2990
rect 123116 2926 123168 2932
rect 123128 480 123156 2926
rect 126440 480 126468 4966
rect 129752 480 129780 4966
rect 131040 4690 131068 38694
rect 131028 4684 131080 4690
rect 131028 4626 131080 4632
rect 131776 3126 131804 38830
rect 131764 3120 131816 3126
rect 131764 3062 131816 3068
rect 131868 3058 131896 38830
rect 136364 6248 136416 6254
rect 136364 6190 136416 6196
rect 133052 3188 133104 3194
rect 133052 3130 133104 3136
rect 131856 3052 131908 3058
rect 131856 2994 131908 3000
rect 133064 480 133092 3130
rect 136376 480 136404 6190
rect 140792 3670 140820 41126
rect 144932 38826 144960 41140
rect 147692 41126 147982 41154
rect 144920 38820 144972 38826
rect 144920 38762 144972 38768
rect 142988 5160 143040 5166
rect 142988 5102 143040 5108
rect 140780 3664 140832 3670
rect 140780 3606 140832 3612
rect 143000 480 143028 5102
rect 146484 3664 146536 3670
rect 146484 3606 146536 3612
rect 146496 480 146524 3606
rect 147692 2990 147720 41126
rect 151004 40662 151032 41140
rect 150992 40656 151044 40662
rect 150992 40598 151044 40604
rect 154132 38826 154160 41140
rect 159928 39982 159956 41140
rect 159916 39976 159968 39982
rect 159916 39918 159968 39924
rect 166000 39681 166028 41140
rect 168760 41138 169142 41154
rect 168748 41132 169142 41138
rect 168800 41126 169142 41132
rect 168748 41074 168800 41080
rect 165986 39672 166042 39681
rect 165986 39607 166042 39616
rect 159364 38956 159416 38962
rect 159364 38898 159416 38904
rect 154120 38820 154172 38826
rect 154120 38762 154172 38768
rect 153108 3596 153160 3602
rect 153108 3538 153160 3544
rect 156420 3596 156472 3602
rect 156420 3538 156472 3544
rect 149796 3256 149848 3262
rect 149796 3198 149848 3204
rect 147680 2984 147732 2990
rect 147680 2926 147732 2932
rect 149808 480 149836 3198
rect 153120 480 153148 3538
rect 156432 480 156460 3538
rect 159376 3262 159404 38898
rect 166356 3392 166408 3398
rect 166356 3334 166408 3340
rect 159732 3324 159784 3330
rect 159732 3266 159784 3272
rect 159364 3256 159416 3262
rect 159364 3198 159416 3204
rect 159744 480 159772 3266
rect 163044 3120 163096 3126
rect 163044 3062 163096 3068
rect 163056 480 163084 3062
rect 166368 480 166396 3334
rect 169680 480 169708 42094
rect 191840 42016 191892 42022
rect 191840 41958 191892 41964
rect 172072 38894 172100 41140
rect 175292 39681 175320 41140
rect 175278 39672 175334 39681
rect 175278 39607 175334 39616
rect 178144 39098 178172 41140
rect 178132 39092 178184 39098
rect 178132 39034 178184 39040
rect 181272 39030 181300 41140
rect 184322 41126 184888 41154
rect 181260 39024 181312 39030
rect 181260 38966 181312 38972
rect 172060 38888 172112 38894
rect 172060 38830 172112 38836
rect 182824 38820 182876 38826
rect 182824 38762 182876 38768
rect 179604 3392 179656 3398
rect 179604 3334 179656 3340
rect 176292 3188 176344 3194
rect 176292 3130 176344 3136
rect 176304 480 176332 3130
rect 179616 480 179644 3334
rect 182836 3126 182864 38762
rect 183100 4140 183152 4146
rect 183100 4082 183152 4088
rect 182824 3120 182876 3126
rect 182824 3062 182876 3068
rect 183112 480 183140 4082
rect 184860 3058 184888 41126
rect 186332 41126 187358 41154
rect 186332 5370 186360 41126
rect 190288 39642 190316 41140
rect 190276 39636 190328 39642
rect 190276 39578 190328 39584
rect 191852 16574 191880 41958
rect 193232 41126 193430 41154
rect 191852 16546 192616 16574
rect 187606 10296 187662 10305
rect 187606 10231 187662 10240
rect 186320 5364 186372 5370
rect 186320 5306 186372 5312
rect 187620 3262 187648 10231
rect 189724 4072 189776 4078
rect 189724 4014 189776 4020
rect 186412 3256 186464 3262
rect 186412 3198 186464 3204
rect 187608 3256 187660 3262
rect 187608 3198 187660 3204
rect 184848 3052 184900 3058
rect 184848 2994 184900 3000
rect 186424 480 186452 3198
rect 189736 480 189764 4014
rect 192588 490 192616 16546
rect 193232 3194 193260 41126
rect 196084 16574 196112 42366
rect 223698 42350 223946 42378
rect 284022 42392 284078 42401
rect 223946 42327 224002 42336
rect 231860 42356 231912 42362
rect 231860 42298 231912 42304
rect 277308 42356 277360 42362
rect 371698 42392 371754 42401
rect 284078 42350 284142 42378
rect 284022 42327 284078 42336
rect 371754 42350 372094 42378
rect 405554 42392 405610 42401
rect 379428 42366 379480 42372
rect 371698 42327 371754 42336
rect 277308 42298 277360 42304
rect 230110 42120 230166 42129
rect 229770 42078 230110 42106
rect 230110 42055 230166 42064
rect 196360 39710 196388 41140
rect 198752 41126 199318 41154
rect 202538 41126 202828 41154
rect 196348 39704 196400 39710
rect 196348 39646 196400 39652
rect 196084 16546 196388 16574
rect 193220 3188 193272 3194
rect 193220 3130 193272 3136
rect 192864 598 193076 626
rect 192864 490 192892 598
rect -10 -960 102 480
rect 3302 -960 3414 480
rect 6614 -960 6726 480
rect 9926 -960 10038 480
rect 13238 -960 13350 480
rect 16550 -960 16662 480
rect 19862 -960 19974 480
rect 23174 -960 23286 480
rect 26486 -960 26598 480
rect 29798 -960 29910 480
rect 33110 -960 33222 480
rect 36606 -960 36718 480
rect 39918 -960 40030 480
rect 43230 -960 43342 480
rect 46542 -960 46654 480
rect 49854 -960 49966 480
rect 53166 -960 53278 480
rect 56478 -960 56590 480
rect 59790 -960 59902 480
rect 63102 -960 63214 480
rect 66414 -960 66526 480
rect 69726 -960 69838 480
rect 73222 -960 73334 480
rect 76534 -960 76646 480
rect 79846 -960 79958 480
rect 83158 -960 83270 480
rect 86470 -960 86582 480
rect 89782 -960 89894 480
rect 93094 -960 93206 480
rect 96406 -960 96518 480
rect 99718 -960 99830 480
rect 103030 -960 103142 480
rect 106342 -960 106454 480
rect 109838 -960 109950 480
rect 113150 -960 113262 480
rect 116462 -960 116574 480
rect 119774 -960 119886 480
rect 123086 -960 123198 480
rect 126398 -960 126510 480
rect 129710 -960 129822 480
rect 133022 -960 133134 480
rect 136334 -960 136446 480
rect 139646 -960 139758 480
rect 142958 -960 143070 480
rect 146454 -960 146566 480
rect 149766 -960 149878 480
rect 153078 -960 153190 480
rect 156390 -960 156502 480
rect 159702 -960 159814 480
rect 163014 -960 163126 480
rect 166326 -960 166438 480
rect 169638 -960 169750 480
rect 172950 -960 173062 480
rect 176262 -960 176374 480
rect 179574 -960 179686 480
rect 183070 -960 183182 480
rect 186382 -960 186494 480
rect 189694 -960 189806 480
rect 192588 462 192892 490
rect 193048 480 193076 598
rect 196360 480 196388 16546
rect 198752 3398 198780 41126
rect 198740 3392 198792 3398
rect 198740 3334 198792 3340
rect 202800 3194 202828 41126
rect 205468 39098 205496 41140
rect 208596 39710 208624 41140
rect 208584 39704 208636 39710
rect 208584 39646 208636 39652
rect 211540 39642 211568 41140
rect 211528 39636 211580 39642
rect 211528 39578 211580 39584
rect 214576 39574 214604 41140
rect 217612 39574 217640 41140
rect 219452 41126 220662 41154
rect 226352 41126 226734 41154
rect 214564 39568 214616 39574
rect 214564 39510 214616 39516
rect 217600 39568 217652 39574
rect 217600 39510 217652 39516
rect 205456 39092 205508 39098
rect 205456 39034 205508 39040
rect 213826 8936 213882 8945
rect 213826 8871 213882 8880
rect 209594 5128 209650 5137
rect 209594 5063 209650 5072
rect 206284 4072 206336 4078
rect 202970 4040 203026 4049
rect 206284 4014 206336 4020
rect 202970 3975 203026 3984
rect 202788 3188 202840 3194
rect 202788 3130 202840 3136
rect 199660 3052 199712 3058
rect 199660 2994 199712 3000
rect 199672 480 199700 2994
rect 202984 480 203012 3975
rect 206296 480 206324 4014
rect 209608 480 209636 5063
rect 213840 2990 213868 8871
rect 219452 4078 219480 41126
rect 226352 41070 226380 41126
rect 226340 41064 226392 41070
rect 226340 41006 226392 41012
rect 231872 16574 231900 42298
rect 275218 41274 275600 41290
rect 275218 41268 275612 41274
rect 275218 41262 275560 41268
rect 275560 41210 275612 41216
rect 232792 41002 232820 41140
rect 234632 41126 235750 41154
rect 232780 40996 232832 41002
rect 232780 40938 232832 40944
rect 231872 16546 232544 16574
rect 229652 5364 229704 5370
rect 229652 5306 229704 5312
rect 219716 4684 219768 4690
rect 219716 4626 219768 4632
rect 226340 4684 226392 4690
rect 226340 4626 226392 4632
rect 219440 4072 219492 4078
rect 219440 4014 219492 4020
rect 213828 2984 213880 2990
rect 213828 2926 213880 2932
rect 216220 2984 216272 2990
rect 216220 2926 216272 2932
rect 216232 480 216260 2926
rect 219728 480 219756 4626
rect 223028 4072 223080 4078
rect 223028 4014 223080 4020
rect 223040 480 223068 4014
rect 226352 480 226380 4626
rect 229664 480 229692 5306
rect 232516 490 232544 16546
rect 234632 4078 234660 41126
rect 238772 41002 238800 41140
rect 238760 40996 238812 41002
rect 238760 40938 238812 40944
rect 241808 39166 241836 41140
rect 244858 41138 245240 41154
rect 244858 41132 245252 41138
rect 244858 41126 245200 41132
rect 245200 41074 245252 41080
rect 247972 39166 248000 41140
rect 250824 39234 250852 41140
rect 250812 39228 250864 39234
rect 250812 39170 250864 39176
rect 241796 39160 241848 39166
rect 241796 39102 241848 39108
rect 247960 39160 248012 39166
rect 247960 39102 248012 39108
rect 254044 38826 254072 41140
rect 256988 39409 257016 41140
rect 256974 39400 257030 39409
rect 256974 39335 257030 39344
rect 260116 39234 260144 41140
rect 263074 41126 263548 41154
rect 260104 39228 260156 39234
rect 260104 39170 260156 39176
rect 259460 39160 259512 39166
rect 259460 39102 259512 39108
rect 254032 38820 254084 38826
rect 254032 38762 254084 38768
rect 255228 38820 255280 38826
rect 255228 38762 255280 38768
rect 246210 6352 246266 6361
rect 246210 6287 246266 6296
rect 242900 5500 242952 5506
rect 242900 5442 242952 5448
rect 239586 5264 239642 5273
rect 239586 5199 239642 5208
rect 234620 4072 234672 4078
rect 234620 4014 234672 4020
rect 236276 4004 236328 4010
rect 236276 3946 236328 3952
rect 232792 598 233004 626
rect 232792 490 232820 598
rect 193006 -960 193118 480
rect 196318 -960 196430 480
rect 199630 -960 199742 480
rect 202942 -960 203054 480
rect 206254 -960 206366 480
rect 209566 -960 209678 480
rect 212878 -960 212990 480
rect 216190 -960 216302 480
rect 219686 -960 219798 480
rect 222998 -960 223110 480
rect 226310 -960 226422 480
rect 229622 -960 229734 480
rect 232516 462 232820 490
rect 232976 480 233004 598
rect 236288 480 236316 3946
rect 239600 480 239628 5199
rect 242912 480 242940 5442
rect 246224 480 246252 6287
rect 255240 4078 255268 38762
rect 259472 16574 259500 39102
rect 259472 16546 259684 16574
rect 256332 4752 256384 4758
rect 256332 4694 256384 4700
rect 255228 4072 255280 4078
rect 249522 4040 249578 4049
rect 255228 4014 255280 4020
rect 249522 3975 249578 3984
rect 249536 480 249564 3975
rect 252836 3936 252888 3942
rect 252836 3878 252888 3884
rect 252848 480 252876 3878
rect 256344 480 256372 4694
rect 259656 480 259684 16546
rect 262956 4140 263008 4146
rect 262956 4082 263008 4088
rect 262968 480 262996 4082
rect 263520 3398 263548 41126
rect 266188 8294 266216 41140
rect 269146 41126 269528 41154
rect 269500 41070 269528 41126
rect 269488 41064 269540 41070
rect 269488 41006 269540 41012
rect 272260 39030 272288 41140
rect 272248 39024 272300 39030
rect 272248 38966 272300 38972
rect 266268 38956 266320 38962
rect 266268 38898 266320 38904
rect 266176 8288 266228 8294
rect 266176 8230 266228 8236
rect 263508 3392 263560 3398
rect 263508 3334 263560 3340
rect 266280 480 266308 38898
rect 269120 19984 269172 19990
rect 269120 19926 269172 19932
rect 269132 490 269160 19926
rect 277320 4010 277348 42298
rect 320180 42288 320232 42294
rect 333888 42288 333940 42294
rect 320232 42236 320574 42242
rect 320180 42230 320574 42236
rect 333888 42230 333940 42236
rect 320192 42214 320574 42230
rect 305920 41336 305972 41342
rect 305578 41284 305920 41290
rect 305578 41278 305972 41284
rect 305578 41262 305960 41278
rect 329196 41200 329248 41206
rect 277412 41126 278070 41154
rect 276204 4004 276256 4010
rect 276204 3946 276256 3952
rect 277308 4004 277360 4010
rect 277308 3946 277360 3952
rect 272892 3936 272944 3942
rect 272892 3878 272944 3884
rect 269408 598 269620 626
rect 269408 490 269436 598
rect 232934 -960 233046 480
rect 236246 -960 236358 480
rect 239558 -960 239670 480
rect 242870 -960 242982 480
rect 246182 -960 246294 480
rect 249494 -960 249606 480
rect 252806 -960 252918 480
rect 256302 -960 256414 480
rect 259614 -960 259726 480
rect 262926 -960 263038 480
rect 266238 -960 266350 480
rect 269132 462 269436 490
rect 269592 480 269620 598
rect 272904 480 272932 3878
rect 276216 480 276244 3946
rect 277412 3942 277440 41126
rect 281276 39166 281304 41140
rect 285678 40624 285734 40633
rect 285678 40559 285734 40568
rect 281264 39160 281316 39166
rect 281264 39102 281316 39108
rect 285692 39098 285720 40559
rect 287348 39545 287376 41140
rect 287334 39536 287390 39545
rect 287334 39471 287390 39480
rect 290292 39098 290320 41140
rect 285680 39092 285732 39098
rect 285680 39034 285732 39040
rect 290280 39092 290332 39098
rect 290280 39034 290332 39040
rect 293328 38962 293356 41140
rect 295444 41126 296286 41154
rect 293316 38956 293368 38962
rect 293316 38898 293368 38904
rect 287702 33552 287758 33561
rect 287702 33487 287758 33496
rect 287716 31074 287744 33487
rect 279424 31068 279476 31074
rect 279424 31010 279476 31016
rect 287704 31068 287756 31074
rect 287704 31010 287756 31016
rect 279436 19990 279464 31010
rect 279424 19984 279476 19990
rect 279424 19926 279476 19932
rect 282828 5500 282880 5506
rect 282828 5442 282880 5448
rect 277400 3936 277452 3942
rect 277400 3878 277452 3884
rect 279516 3936 279568 3942
rect 279516 3878 279568 3884
rect 279528 480 279556 3878
rect 282840 480 282868 5442
rect 284300 4616 284352 4622
rect 284300 4558 284352 4564
rect 284312 3058 284340 4558
rect 286140 4004 286192 4010
rect 286140 3946 286192 3952
rect 284300 3052 284352 3058
rect 284300 2994 284352 3000
rect 286152 480 286180 3946
rect 295444 3330 295472 41126
rect 296260 4752 296312 4758
rect 296260 4694 296312 4700
rect 289452 3324 289504 3330
rect 289452 3266 289504 3272
rect 292948 3324 293000 3330
rect 292948 3266 293000 3272
rect 295432 3324 295484 3330
rect 295432 3266 295484 3272
rect 289464 480 289492 3266
rect 292960 480 292988 3266
rect 296272 480 296300 4694
rect 299492 4690 299520 41140
rect 302344 39302 302372 41140
rect 308508 39953 308536 41140
rect 311650 41126 311848 41154
rect 308494 39944 308550 39953
rect 308494 39879 308550 39888
rect 302332 39296 302384 39302
rect 302332 39238 302384 39244
rect 301504 39024 301556 39030
rect 301504 38966 301556 38972
rect 299480 4684 299532 4690
rect 299480 4626 299532 4632
rect 299572 4684 299624 4690
rect 299572 4626 299624 4632
rect 299584 480 299612 4626
rect 301516 3058 301544 38966
rect 309506 6488 309562 6497
rect 309506 6423 309562 6432
rect 302882 5536 302938 5545
rect 302882 5471 302938 5480
rect 301504 3052 301556 3058
rect 301504 2994 301556 3000
rect 302896 480 302924 5471
rect 306196 3120 306248 3126
rect 306196 3062 306248 3068
rect 306208 480 306236 3062
rect 309520 480 309548 6423
rect 311820 3126 311848 41126
rect 314580 39982 314608 41140
rect 314568 39976 314620 39982
rect 314568 39918 314620 39924
rect 316040 39976 316092 39982
rect 316040 39918 316092 39924
rect 316052 16574 316080 39918
rect 317524 39273 317552 41140
rect 323610 41126 324268 41154
rect 326738 41126 327028 41154
rect 329248 41148 329590 41154
rect 329196 41142 329590 41148
rect 329208 41126 329590 41142
rect 317510 39264 317566 39273
rect 317510 39199 317566 39208
rect 320824 22092 320876 22098
rect 320824 22034 320876 22040
rect 316052 16546 316172 16574
rect 312820 3324 312872 3330
rect 312820 3266 312872 3272
rect 311808 3120 311860 3126
rect 311808 3062 311860 3068
rect 312832 480 312860 3266
rect 316144 480 316172 16546
rect 320836 4690 320864 22034
rect 320824 4684 320876 4690
rect 320824 4626 320876 4632
rect 324240 3874 324268 41126
rect 326620 23588 326672 23594
rect 326620 23530 326672 23536
rect 326632 22166 326660 23530
rect 326620 22160 326672 22166
rect 326620 22102 326672 22108
rect 326344 15156 326396 15162
rect 326344 15098 326396 15104
rect 326356 4622 326384 15098
rect 326344 4616 326396 4622
rect 326344 4558 326396 4564
rect 319444 3868 319496 3874
rect 319444 3810 319496 3816
rect 324228 3868 324280 3874
rect 324228 3810 324280 3816
rect 326068 3868 326120 3874
rect 326068 3810 326120 3816
rect 319456 480 319484 3810
rect 322756 3732 322808 3738
rect 322756 3674 322808 3680
rect 322768 480 322796 3674
rect 326080 480 326108 3810
rect 327000 3738 327028 41126
rect 332796 39302 332824 41140
rect 332784 39296 332836 39302
rect 332784 39238 332836 39244
rect 332600 27668 332652 27674
rect 332600 27610 332652 27616
rect 331220 25356 331272 25362
rect 331220 25298 331272 25304
rect 331232 23594 331260 25298
rect 331220 23588 331272 23594
rect 331220 23530 331272 23536
rect 332612 23526 332640 27610
rect 329840 23520 329892 23526
rect 329840 23462 329892 23468
rect 332600 23520 332652 23526
rect 332600 23462 332652 23468
rect 329852 19258 329880 23462
rect 329484 19230 329880 19258
rect 329484 15230 329512 19230
rect 329472 15224 329524 15230
rect 329472 15166 329524 15172
rect 333900 3738 333928 42230
rect 348238 41440 348294 41449
rect 348238 41375 348294 41384
rect 335648 39438 335676 41140
rect 338776 39506 338804 41140
rect 340892 41126 341734 41154
rect 338764 39500 338816 39506
rect 338764 39442 338816 39448
rect 335636 39432 335688 39438
rect 335636 39374 335688 39380
rect 340512 34468 340564 34474
rect 340512 34410 340564 34416
rect 340524 31822 340552 34410
rect 340512 31816 340564 31822
rect 340512 31758 340564 31764
rect 336004 31748 336056 31754
rect 336004 31690 336056 31696
rect 339684 31748 339736 31754
rect 339684 31690 339736 31696
rect 336016 25362 336044 31690
rect 339696 29850 339724 31690
rect 338028 29844 338080 29850
rect 338028 29786 338080 29792
rect 339684 29844 339736 29850
rect 339684 29786 339736 29792
rect 338040 27674 338068 29786
rect 338028 27668 338080 27674
rect 338028 27610 338080 27616
rect 336004 25356 336056 25362
rect 336004 25298 336056 25304
rect 340144 15224 340196 15230
rect 340144 15166 340196 15172
rect 340156 4758 340184 15166
rect 340144 4752 340196 4758
rect 340144 4694 340196 4700
rect 339498 3904 339554 3913
rect 339498 3839 339554 3848
rect 326988 3732 327040 3738
rect 326988 3674 327040 3680
rect 329564 3732 329616 3738
rect 329564 3674 329616 3680
rect 332876 3732 332928 3738
rect 332876 3674 332928 3680
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 336188 3732 336240 3738
rect 336188 3674 336240 3680
rect 329576 480 329604 3674
rect 332888 480 332916 3674
rect 336200 480 336228 3674
rect 339512 480 339540 3839
rect 340892 3806 340920 41126
rect 344940 39506 344968 41140
rect 347792 40934 347820 41140
rect 347780 40928 347832 40934
rect 347780 40870 347832 40876
rect 348252 40050 348280 41375
rect 366456 41200 366508 41206
rect 351012 40934 351040 41140
rect 351000 40928 351052 40934
rect 351000 40870 351052 40876
rect 353864 40361 353892 41140
rect 356914 41126 357388 41154
rect 360042 41126 360148 41154
rect 366114 41148 366456 41154
rect 366114 41142 366508 41148
rect 353850 40352 353906 40361
rect 353850 40287 353906 40296
rect 354954 40352 355010 40361
rect 354954 40287 355010 40296
rect 354968 40050 354996 40287
rect 345664 40044 345716 40050
rect 345664 39986 345716 39992
rect 348240 40044 348292 40050
rect 348240 39986 348292 39992
rect 352380 40044 352432 40050
rect 352380 39986 352432 39992
rect 354956 40044 355008 40050
rect 354956 39986 355008 39992
rect 344928 39500 344980 39506
rect 344928 39442 344980 39448
rect 343548 35964 343600 35970
rect 343548 35906 343600 35912
rect 343560 33182 343588 35906
rect 343640 35284 343692 35290
rect 343640 35226 343692 35232
rect 341524 33176 341576 33182
rect 341524 33118 341576 33124
rect 343548 33176 343600 33182
rect 343548 33118 343600 33124
rect 341536 15230 341564 33118
rect 343652 31822 343680 35226
rect 345676 34542 345704 39986
rect 350538 39128 350594 39137
rect 350538 39063 350594 39072
rect 350552 38350 350580 39063
rect 346308 38344 346360 38350
rect 346308 38286 346360 38292
rect 350540 38344 350592 38350
rect 350540 38286 350592 38292
rect 346320 35970 346348 38286
rect 352392 37942 352420 39986
rect 349988 37936 350040 37942
rect 349988 37878 350040 37884
rect 352380 37936 352432 37942
rect 352380 37878 352432 37884
rect 346308 35964 346360 35970
rect 346308 35906 346360 35912
rect 350000 35290 350028 37878
rect 354586 35864 354642 35873
rect 354586 35799 354642 35808
rect 349988 35284 350040 35290
rect 349988 35226 350040 35232
rect 349160 35216 349212 35222
rect 349160 35158 349212 35164
rect 345664 34536 345716 34542
rect 345664 34478 345716 34484
rect 343640 31816 343692 31822
rect 343640 31758 343692 31764
rect 349172 16574 349200 35158
rect 354600 26353 354628 35799
rect 354586 26344 354642 26353
rect 354586 26279 354642 26288
rect 354586 26208 354642 26217
rect 354586 26143 354642 26152
rect 354600 16697 354628 26143
rect 354586 16688 354642 16697
rect 354586 16623 354642 16632
rect 349172 16546 349476 16574
rect 341524 15224 341576 15230
rect 341524 15166 341576 15172
rect 340880 3800 340932 3806
rect 340880 3742 340932 3748
rect 342812 3256 342864 3262
rect 342812 3198 342864 3204
rect 342824 480 342852 3198
rect 346124 3188 346176 3194
rect 346124 3130 346176 3136
rect 346136 480 346164 3130
rect 349448 480 349476 16546
rect 354586 16552 354642 16561
rect 354586 16487 354642 16496
rect 354600 7041 354628 16487
rect 354586 7032 354642 7041
rect 354586 6967 354642 6976
rect 352748 5432 352800 5438
rect 352748 5374 352800 5380
rect 356060 5432 356112 5438
rect 356060 5374 356112 5380
rect 352760 480 352788 5374
rect 356072 480 356100 5374
rect 357360 4690 357388 41126
rect 357348 4684 357400 4690
rect 357348 4626 357400 4632
rect 359370 3904 359426 3913
rect 359370 3839 359426 3848
rect 359384 480 359412 3839
rect 360120 3262 360148 41126
rect 362972 39030 363000 41140
rect 366114 41126 366496 41142
rect 369044 39438 369072 41140
rect 369032 39432 369084 39438
rect 369032 39374 369084 39380
rect 375116 39302 375144 41140
rect 367744 39296 367796 39302
rect 367744 39238 367796 39244
rect 375104 39296 375156 39302
rect 375104 39238 375156 39244
rect 362960 39024 363012 39030
rect 362960 38966 363012 38972
rect 367756 3806 367784 39238
rect 372620 39024 372672 39030
rect 372620 38966 372672 38972
rect 368480 36576 368532 36582
rect 368480 36518 368532 36524
rect 368492 16574 368520 36518
rect 372632 16574 372660 38966
rect 378152 38729 378180 41140
rect 378138 38720 378194 38729
rect 378138 38655 378194 38664
rect 368492 16546 369072 16574
rect 372632 16546 372844 16574
rect 367744 3800 367796 3806
rect 367744 3742 367796 3748
rect 360108 3256 360160 3262
rect 360108 3198 360160 3204
rect 366180 3256 366232 3262
rect 366180 3198 366232 3204
rect 362682 3088 362738 3097
rect 362682 3023 362738 3032
rect 362696 480 362724 3023
rect 366192 480 366220 3198
rect 369044 490 369072 16546
rect 369320 598 369532 626
rect 369320 490 369348 598
rect 269550 -960 269662 480
rect 272862 -960 272974 480
rect 276174 -960 276286 480
rect 279486 -960 279598 480
rect 282798 -960 282910 480
rect 286110 -960 286222 480
rect 289422 -960 289534 480
rect 292918 -960 293030 480
rect 296230 -960 296342 480
rect 299542 -960 299654 480
rect 302854 -960 302966 480
rect 306166 -960 306278 480
rect 309478 -960 309590 480
rect 312790 -960 312902 480
rect 316102 -960 316214 480
rect 319414 -960 319526 480
rect 322726 -960 322838 480
rect 326038 -960 326150 480
rect 329534 -960 329646 480
rect 332846 -960 332958 480
rect 336158 -960 336270 480
rect 339470 -960 339582 480
rect 342782 -960 342894 480
rect 346094 -960 346206 480
rect 349406 -960 349518 480
rect 352718 -960 352830 480
rect 356030 -960 356142 480
rect 359342 -960 359454 480
rect 362654 -960 362766 480
rect 366150 -960 366262 480
rect 369044 462 369348 490
rect 369504 480 369532 598
rect 372816 480 372844 16546
rect 376116 6316 376168 6322
rect 376116 6258 376168 6264
rect 376128 480 376156 6258
rect 379440 480 379468 42366
rect 405490 42350 405554 42378
rect 405554 42327 405610 42336
rect 382280 42220 382332 42226
rect 382280 42162 382332 42168
rect 395988 42220 396040 42226
rect 395988 42162 396040 42168
rect 381096 40225 381124 41140
rect 381082 40216 381138 40225
rect 381082 40151 381138 40160
rect 382292 490 382320 42162
rect 384330 41410 384712 41426
rect 384330 41404 384724 41410
rect 384330 41398 384672 41404
rect 384672 41346 384724 41352
rect 387260 39302 387288 41140
rect 390296 40089 390324 41140
rect 393332 40089 393360 41140
rect 390282 40080 390338 40089
rect 390282 40015 390338 40024
rect 393318 40080 393374 40089
rect 393318 40015 393374 40024
rect 385040 39296 385092 39302
rect 385040 39238 385092 39244
rect 387248 39296 387300 39302
rect 387248 39238 387300 39244
rect 385052 16574 385080 39238
rect 385052 16546 385632 16574
rect 382568 598 382780 626
rect 382568 490 382596 598
rect 369462 -960 369574 480
rect 372774 -960 372886 480
rect 376086 -960 376198 480
rect 379398 -960 379510 480
rect 382292 462 382596 490
rect 382752 480 382780 598
rect 385604 490 385632 16546
rect 389364 4752 389416 4758
rect 389364 4694 389416 4700
rect 385880 598 386092 626
rect 385880 490 385908 598
rect 382710 -960 382822 480
rect 385604 462 385908 490
rect 386064 480 386092 598
rect 389376 480 389404 4694
rect 392674 2952 392730 2961
rect 392674 2887 392730 2896
rect 392688 480 392716 2887
rect 396000 480 396028 42162
rect 436008 42016 436060 42022
rect 436008 41958 436060 41964
rect 509148 42016 509200 42022
rect 509148 41958 509200 41964
rect 536748 42016 536800 42022
rect 536748 41958 536800 41964
rect 396092 41126 396198 41154
rect 399418 41126 400168 41154
rect 402362 41126 402928 41154
rect 396092 5302 396120 41126
rect 396080 5296 396132 5302
rect 396080 5238 396132 5244
rect 400140 3874 400168 41126
rect 400128 3868 400180 3874
rect 400128 3810 400180 3816
rect 402900 3262 402928 41126
rect 408328 40866 408356 41140
rect 408316 40860 408368 40866
rect 408316 40802 408368 40808
rect 411456 40798 411484 41140
rect 411444 40792 411496 40798
rect 411444 40734 411496 40740
rect 414492 38826 414520 41140
rect 417528 39846 417556 41140
rect 420472 40730 420500 41140
rect 420460 40724 420512 40730
rect 420460 40666 420512 40672
rect 417516 39840 417568 39846
rect 417516 39782 417568 39788
rect 423692 39137 423720 41140
rect 426636 39846 426664 41140
rect 429672 39914 429700 41140
rect 429660 39908 429712 39914
rect 429660 39850 429712 39856
rect 426624 39840 426676 39846
rect 426624 39782 426676 39788
rect 423678 39128 423734 39137
rect 423678 39063 423734 39072
rect 432616 38865 432644 41140
rect 435652 39030 435680 41140
rect 435640 39024 435692 39030
rect 435640 38966 435692 38972
rect 432602 38856 432658 38865
rect 414480 38820 414532 38826
rect 414480 38762 414532 38768
rect 415308 38820 415360 38826
rect 432602 38791 432658 38800
rect 415308 38762 415360 38768
rect 406108 5296 406160 5302
rect 406108 5238 406160 5244
rect 402888 3256 402940 3262
rect 402888 3198 402940 3204
rect 399300 3120 399352 3126
rect 399300 3062 399352 3068
rect 399312 480 399340 3062
rect 402794 2952 402850 2961
rect 402794 2887 402850 2896
rect 402808 480 402836 2887
rect 406120 480 406148 5238
rect 409420 5228 409472 5234
rect 409420 5170 409472 5176
rect 409432 480 409460 5170
rect 415320 3194 415348 38762
rect 436020 6914 436048 41958
rect 438780 33114 438808 41140
rect 441632 40594 441660 41140
rect 441620 40588 441672 40594
rect 441620 40530 441672 40536
rect 439504 39840 439556 39846
rect 439504 39782 439556 39788
rect 438768 33108 438820 33114
rect 438768 33050 438820 33056
rect 435928 6886 436048 6914
rect 419354 4992 419410 5001
rect 419354 4927 419410 4936
rect 415308 3188 415360 3194
rect 415308 3130 415360 3136
rect 412730 3088 412786 3097
rect 412730 3023 412786 3032
rect 416044 3052 416096 3058
rect 412744 480 412772 3023
rect 416044 2994 416096 3000
rect 416056 480 416084 2994
rect 419368 480 419396 4927
rect 429292 3188 429344 3194
rect 429292 3130 429344 3136
rect 425978 3088 426034 3097
rect 425978 3023 426034 3032
rect 425992 480 426020 3023
rect 429304 480 429332 3130
rect 432602 3088 432658 3097
rect 432602 3023 432658 3032
rect 432616 480 432644 3023
rect 435928 480 435956 6886
rect 439410 3224 439466 3233
rect 439516 3194 439544 39782
rect 443644 39364 443696 39370
rect 443644 39306 443696 39312
rect 442724 4684 442776 4690
rect 442724 4626 442776 4632
rect 439410 3159 439466 3168
rect 439504 3188 439556 3194
rect 439424 480 439452 3159
rect 439504 3130 439556 3136
rect 442736 480 442764 4626
rect 443656 3126 443684 39306
rect 444852 38894 444880 41140
rect 447810 41126 448468 41154
rect 444840 38888 444892 38894
rect 444840 38830 444892 38836
rect 446036 3188 446088 3194
rect 446036 3130 446088 3136
rect 443644 3120 443696 3126
rect 443644 3062 443696 3068
rect 446048 480 446076 3130
rect 448440 3058 448468 41126
rect 450924 39846 450952 41140
rect 450912 39840 450964 39846
rect 450912 39782 450964 39788
rect 453776 39778 453804 41140
rect 456812 41126 456918 41154
rect 453764 39772 453816 39778
rect 453764 39714 453816 39720
rect 451924 39024 451976 39030
rect 451924 38966 451976 38972
rect 449808 37936 449860 37942
rect 449808 37878 449860 37884
rect 449820 3194 449848 37878
rect 451936 3194 451964 38966
rect 456812 6254 456840 41126
rect 459940 39778 459968 41140
rect 459928 39772 459980 39778
rect 459928 39714 459980 39720
rect 462976 39409 463004 41140
rect 465920 40390 465948 41140
rect 469140 40390 469168 41140
rect 465908 40384 465960 40390
rect 465908 40326 465960 40332
rect 469128 40384 469180 40390
rect 469128 40326 469180 40332
rect 462962 39400 463018 39409
rect 462962 39335 463018 39344
rect 471992 39001 472020 41140
rect 474936 40322 474964 41140
rect 477512 41126 478078 41154
rect 480272 41126 481022 41154
rect 474924 40316 474976 40322
rect 474924 40258 474976 40264
rect 471978 38992 472034 39001
rect 471978 38927 472034 38936
rect 456800 6248 456852 6254
rect 456800 6190 456852 6196
rect 452660 5092 452712 5098
rect 452660 5034 452712 5040
rect 449348 3188 449400 3194
rect 449348 3130 449400 3136
rect 449808 3188 449860 3194
rect 449808 3130 449860 3136
rect 451924 3188 451976 3194
rect 451924 3130 451976 3136
rect 448428 3052 448480 3058
rect 448428 2994 448480 3000
rect 449360 480 449388 3130
rect 452672 480 452700 5034
rect 476026 4992 476082 5001
rect 476026 4927 476082 4936
rect 469220 3528 469272 3534
rect 469220 3470 469272 3476
rect 465908 3256 465960 3262
rect 465908 3198 465960 3204
rect 455972 3188 456024 3194
rect 455972 3130 456024 3136
rect 462596 3188 462648 3194
rect 462596 3130 462648 3136
rect 455984 480 456012 3130
rect 459282 3088 459338 3097
rect 459282 3023 459338 3032
rect 459296 480 459324 3023
rect 462608 480 462636 3130
rect 465920 480 465948 3198
rect 469232 480 469260 3470
rect 472532 3052 472584 3058
rect 472532 2994 472584 3000
rect 472544 480 472572 2994
rect 476040 480 476068 4927
rect 477512 3670 477540 41126
rect 480272 4962 480300 41126
rect 484136 38826 484164 41140
rect 482928 38820 482980 38826
rect 482928 38762 482980 38768
rect 484124 38820 484176 38826
rect 484124 38762 484176 38768
rect 482940 6914 482968 38762
rect 482664 6886 482968 6914
rect 480260 4956 480312 4962
rect 480260 4898 480312 4904
rect 477500 3664 477552 3670
rect 477500 3606 477552 3612
rect 479338 3360 479394 3369
rect 479338 3295 479394 3304
rect 479352 480 479380 3295
rect 482664 480 482692 6886
rect 487172 4146 487200 41140
rect 490300 39030 490328 41140
rect 493244 40594 493272 41140
rect 493232 40588 493284 40594
rect 493232 40530 493284 40536
rect 496372 40322 496400 41140
rect 496360 40316 496412 40322
rect 496360 40258 496412 40264
rect 499224 40254 499252 41140
rect 499212 40248 499264 40254
rect 499212 40190 499264 40196
rect 490288 39024 490340 39030
rect 490288 38966 490340 38972
rect 502444 38962 502472 41140
rect 505112 41126 505310 41154
rect 502432 38956 502484 38962
rect 502432 38898 502484 38904
rect 488538 33824 488594 33833
rect 488538 33759 488594 33768
rect 488552 16574 488580 33759
rect 498200 25560 498252 25566
rect 498200 25502 498252 25508
rect 498212 16574 498240 25502
rect 488552 16546 488856 16574
rect 498212 16546 498792 16574
rect 487160 4140 487212 4146
rect 487160 4082 487212 4088
rect 485964 3392 486016 3398
rect 485964 3334 486016 3340
rect 485976 480 486004 3334
rect 488828 490 488856 16546
rect 492588 4072 492640 4078
rect 492588 4014 492640 4020
rect 489104 598 489316 626
rect 489104 490 489132 598
rect 386022 -960 386134 480
rect 389334 -960 389446 480
rect 392646 -960 392758 480
rect 395958 -960 396070 480
rect 399270 -960 399382 480
rect 402766 -960 402878 480
rect 406078 -960 406190 480
rect 409390 -960 409502 480
rect 412702 -960 412814 480
rect 416014 -960 416126 480
rect 419326 -960 419438 480
rect 422638 -960 422750 480
rect 425950 -960 426062 480
rect 429262 -960 429374 480
rect 432574 -960 432686 480
rect 435886 -960 435998 480
rect 439382 -960 439494 480
rect 442694 -960 442806 480
rect 446006 -960 446118 480
rect 449318 -960 449430 480
rect 452630 -960 452742 480
rect 455942 -960 456054 480
rect 459254 -960 459366 480
rect 462566 -960 462678 480
rect 465878 -960 465990 480
rect 469190 -960 469302 480
rect 472502 -960 472614 480
rect 475998 -960 476110 480
rect 479310 -960 479422 480
rect 482622 -960 482734 480
rect 485934 -960 486046 480
rect 488828 462 489132 490
rect 489288 480 489316 598
rect 492600 480 492628 4014
rect 495900 3528 495952 3534
rect 495900 3470 495952 3476
rect 495912 480 495940 3470
rect 498764 490 498792 16546
rect 505112 4758 505140 41126
rect 508424 40186 508452 41140
rect 508412 40180 508464 40186
rect 508412 40122 508464 40128
rect 505100 4752 505152 4758
rect 505100 4694 505152 4700
rect 505836 3664 505888 3670
rect 505836 3606 505888 3612
rect 502524 3120 502576 3126
rect 502524 3062 502576 3068
rect 499040 598 499252 626
rect 499040 490 499068 598
rect 489246 -960 489358 480
rect 492558 -960 492670 480
rect 495870 -960 495982 480
rect 498764 462 499068 490
rect 499224 480 499252 598
rect 502536 480 502564 3062
rect 505848 480 505876 3606
rect 509160 480 509188 41958
rect 511460 40050 511488 41140
rect 513288 40724 513340 40730
rect 513288 40666 513340 40672
rect 511448 40044 511500 40050
rect 511448 39986 511500 39992
rect 513300 3058 513328 40666
rect 514404 39370 514432 41140
rect 514392 39364 514444 39370
rect 514392 39306 514444 39312
rect 515954 3632 516010 3641
rect 515954 3567 516010 3576
rect 512644 3052 512696 3058
rect 512644 2994 512696 3000
rect 513288 3052 513340 3058
rect 513288 2994 513340 3000
rect 512656 480 512684 2994
rect 515968 480 515996 3567
rect 517532 3330 517560 41140
rect 520384 40118 520412 41140
rect 523052 41126 523526 41154
rect 526562 41126 527128 41154
rect 520372 40112 520424 40118
rect 520372 40054 520424 40060
rect 519266 3904 519322 3913
rect 519266 3839 519322 3848
rect 517520 3324 517572 3330
rect 517520 3266 517572 3272
rect 519280 480 519308 3839
rect 522580 3460 522632 3466
rect 522580 3402 522632 3408
rect 522592 480 522620 3402
rect 523052 3194 523080 41126
rect 527100 3398 527128 41126
rect 529676 39982 529704 41140
rect 529664 39976 529716 39982
rect 529664 39918 529716 39924
rect 528558 33824 528614 33833
rect 528558 33759 528614 33768
rect 528572 16574 528600 33759
rect 528572 16546 528784 16574
rect 527088 3392 527140 3398
rect 527088 3334 527140 3340
rect 525892 3324 525944 3330
rect 525892 3266 525944 3272
rect 523040 3188 523092 3194
rect 523040 3130 523092 3136
rect 525904 480 525932 3266
rect 528756 490 528784 16546
rect 532620 4078 532648 41140
rect 535748 39914 535776 41140
rect 535736 39908 535788 39914
rect 535736 39850 535788 39856
rect 532608 4072 532660 4078
rect 532608 4014 532660 4020
rect 536760 3466 536788 41958
rect 538312 41472 538364 41478
rect 538312 41414 538364 41420
rect 538324 16574 538352 41414
rect 538692 38826 538720 41140
rect 541820 38894 541848 41140
rect 541808 38888 541860 38894
rect 541808 38830 541860 38836
rect 538680 38820 538732 38826
rect 538680 38762 538732 38768
rect 539508 38820 539560 38826
rect 539508 38762 539560 38768
rect 538324 16546 538720 16574
rect 535828 3460 535880 3466
rect 535828 3402 535880 3408
rect 536748 3460 536800 3466
rect 536748 3402 536800 3408
rect 532516 3256 532568 3262
rect 532516 3198 532568 3204
rect 529032 598 529244 626
rect 529032 490 529060 598
rect 499182 -960 499294 480
rect 502494 -960 502606 480
rect 505806 -960 505918 480
rect 509118 -960 509230 480
rect 512614 -960 512726 480
rect 515926 -960 516038 480
rect 519238 -960 519350 480
rect 522550 -960 522662 480
rect 525862 -960 525974 480
rect 528756 462 529060 490
rect 529216 480 529244 598
rect 532528 480 532556 3198
rect 535840 480 535868 3402
rect 538692 490 538720 16546
rect 539520 4146 539548 38762
rect 542004 4894 542032 143919
rect 542174 117328 542230 117337
rect 542174 117263 542230 117272
rect 542082 95160 542138 95169
rect 542082 95095 542138 95104
rect 542096 6186 542124 95095
rect 542188 44266 542216 117263
rect 542268 73228 542320 73234
rect 542268 73170 542320 73176
rect 542176 44260 542228 44266
rect 542176 44202 542228 44208
rect 542176 43988 542228 43994
rect 542176 43930 542228 43936
rect 542188 43110 542216 43930
rect 542280 43246 542308 73170
rect 542268 43240 542320 43246
rect 542268 43182 542320 43188
rect 542176 43104 542228 43110
rect 542176 43046 542228 43052
rect 542372 41478 542400 664770
rect 542452 663808 542504 663814
rect 542452 663750 542504 663756
rect 542464 42430 542492 663750
rect 542728 663672 542780 663678
rect 542728 663614 542780 663620
rect 542636 662244 542688 662250
rect 542636 662186 542688 662192
rect 542544 660612 542596 660618
rect 542544 660554 542596 660560
rect 542556 660521 542584 660554
rect 542542 660512 542598 660521
rect 542542 660447 542598 660456
rect 542544 660272 542596 660278
rect 542544 660214 542596 660220
rect 542556 530097 542584 660214
rect 542648 633457 542676 662186
rect 542740 660278 542768 663614
rect 542728 660272 542780 660278
rect 542728 660214 542780 660220
rect 542728 659660 542780 659666
rect 542728 659602 542780 659608
rect 542740 641889 542768 659602
rect 542726 641880 542782 641889
rect 542726 641815 542782 641824
rect 542634 633448 542690 633457
rect 542634 633383 542690 633392
rect 542636 620356 542688 620362
rect 542636 620298 542688 620304
rect 542648 615233 542676 620298
rect 542634 615224 542690 615233
rect 542634 615159 542690 615168
rect 542542 530088 542598 530097
rect 542542 530023 542598 530032
rect 542542 524512 542598 524521
rect 542542 524447 542598 524456
rect 542452 42424 542504 42430
rect 542452 42366 542504 42372
rect 542360 41472 542412 41478
rect 542360 41414 542412 41420
rect 542268 38888 542320 38894
rect 542268 38830 542320 38836
rect 542084 6180 542136 6186
rect 542084 6122 542136 6128
rect 541992 4888 542044 4894
rect 541992 4830 542044 4836
rect 539508 4140 539560 4146
rect 539508 4082 539560 4088
rect 542280 4078 542308 38830
rect 542452 4820 542504 4826
rect 542452 4762 542504 4768
rect 542268 4072 542320 4078
rect 542268 4014 542320 4020
rect 538968 598 539180 626
rect 538968 490 538996 598
rect 529174 -960 529286 480
rect 532486 -960 532598 480
rect 535798 -960 535910 480
rect 538692 462 538996 490
rect 539152 480 539180 598
rect 542464 480 542492 4762
rect 542556 4010 542584 524447
rect 542636 505980 542688 505986
rect 542636 505922 542688 505928
rect 542648 503441 542676 505922
rect 542634 503432 542690 503441
rect 542634 503367 542690 503376
rect 542726 484528 542782 484537
rect 542726 484463 542782 484472
rect 542634 480312 542690 480321
rect 542634 480247 542690 480256
rect 542544 4004 542596 4010
rect 542544 3946 542596 3952
rect 542648 3670 542676 480247
rect 542740 43722 542768 484463
rect 542832 301889 542860 700470
rect 542912 700120 542964 700126
rect 542912 700062 542964 700068
rect 542924 350305 542952 700062
rect 543372 663536 543424 663542
rect 543372 663478 543424 663484
rect 543280 661632 543332 661638
rect 543280 661574 543332 661580
rect 543096 661496 543148 661502
rect 543096 661438 543148 661444
rect 543004 661428 543056 661434
rect 543004 661370 543056 661376
rect 542910 350296 542966 350305
rect 542910 350231 542966 350240
rect 543016 336734 543044 661370
rect 543108 355201 543136 661438
rect 543188 660204 543240 660210
rect 543188 660146 543240 660152
rect 543200 382634 543228 660146
rect 543292 422385 543320 661574
rect 543384 659666 543412 663478
rect 543464 662516 543516 662522
rect 543464 662458 543516 662464
rect 543476 660278 543504 662458
rect 543556 660680 543608 660686
rect 543556 660622 543608 660628
rect 543464 660272 543516 660278
rect 543464 660214 543516 660220
rect 543464 660136 543516 660142
rect 543464 660078 543516 660084
rect 543372 659660 543424 659666
rect 543372 659602 543424 659608
rect 543372 659524 543424 659530
rect 543372 659466 543424 659472
rect 543384 485858 543412 659466
rect 543476 547194 543504 660078
rect 543568 600982 543596 660622
rect 543660 655518 543688 700538
rect 543648 655512 543700 655518
rect 543648 655454 543700 655460
rect 543648 651296 543700 651302
rect 543648 651238 543700 651244
rect 543660 651137 543688 651238
rect 543646 651128 543702 651137
rect 543646 651063 543702 651072
rect 543556 600976 543608 600982
rect 543556 600918 543608 600924
rect 543648 597032 543700 597038
rect 543646 597000 543648 597009
rect 543700 597000 543702 597009
rect 543646 596935 543702 596944
rect 543464 547188 543516 547194
rect 543464 547130 543516 547136
rect 543464 543244 543516 543250
rect 543464 543186 543516 543192
rect 543372 485852 543424 485858
rect 543372 485794 543424 485800
rect 543476 458862 543504 543186
rect 543464 458856 543516 458862
rect 543464 458798 543516 458804
rect 543278 422376 543334 422385
rect 543278 422311 543334 422320
rect 543188 382628 543240 382634
rect 543188 382570 543240 382576
rect 543094 355192 543150 355201
rect 543094 355127 543150 355136
rect 543004 336728 543056 336734
rect 543004 336670 543056 336676
rect 542910 305280 542966 305289
rect 542910 305215 542966 305224
rect 542818 301880 542874 301889
rect 542818 301815 542874 301824
rect 542818 291680 542874 291689
rect 542818 291615 542874 291624
rect 542832 44674 542860 291615
rect 542820 44668 542872 44674
rect 542820 44610 542872 44616
rect 542820 44260 542872 44266
rect 542820 44202 542872 44208
rect 542728 43716 542780 43722
rect 542728 43658 542780 43664
rect 542728 43580 542780 43586
rect 542728 43522 542780 43528
rect 542740 40730 542768 43522
rect 542832 43314 542860 44202
rect 542820 43308 542872 43314
rect 542820 43250 542872 43256
rect 542728 40724 542780 40730
rect 542728 40666 542780 40672
rect 542924 5370 542952 305215
rect 543002 202192 543058 202201
rect 543002 202127 543058 202136
rect 542912 5364 542964 5370
rect 542912 5306 542964 5312
rect 542636 3664 542688 3670
rect 542636 3606 542688 3612
rect 543016 3330 543044 202127
rect 543094 198384 543150 198393
rect 543094 198319 543150 198328
rect 543108 3942 543136 198319
rect 543278 153504 543334 153513
rect 543278 153439 543334 153448
rect 543186 140176 543242 140185
rect 543186 140111 543242 140120
rect 543096 3936 543148 3942
rect 543096 3878 543148 3884
rect 543200 3738 543228 140111
rect 543292 42566 543320 153439
rect 543752 109041 543780 700606
rect 543844 252113 543872 700742
rect 543936 458289 543964 700878
rect 544200 700324 544252 700330
rect 544200 700266 544252 700272
rect 544016 663128 544068 663134
rect 544016 663070 544068 663076
rect 544028 660142 544056 663070
rect 544108 662448 544160 662454
rect 544108 662390 544160 662396
rect 544016 660136 544068 660142
rect 544016 660078 544068 660084
rect 544016 659864 544068 659870
rect 544016 659806 544068 659812
rect 544028 655217 544056 659806
rect 544120 659326 544148 662390
rect 544108 659320 544160 659326
rect 544108 659262 544160 659268
rect 544108 659184 544160 659190
rect 544108 659126 544160 659132
rect 544120 655654 544148 659126
rect 544108 655648 544160 655654
rect 544108 655590 544160 655596
rect 544108 655512 544160 655518
rect 544108 655454 544160 655460
rect 544014 655208 544070 655217
rect 544014 655143 544070 655152
rect 544016 655104 544068 655110
rect 544016 655046 544068 655052
rect 543922 458280 543978 458289
rect 543922 458215 543978 458224
rect 543924 435736 543976 435742
rect 543922 435704 543924 435713
rect 543976 435704 543978 435713
rect 543922 435639 543978 435648
rect 543924 431384 543976 431390
rect 543922 431352 543924 431361
rect 543976 431352 543978 431361
rect 543922 431287 543978 431296
rect 544028 426737 544056 655046
rect 544120 630018 544148 655454
rect 544108 630012 544160 630018
rect 544108 629954 544160 629960
rect 544106 628144 544162 628153
rect 544106 628079 544162 628088
rect 544014 426728 544070 426737
rect 544014 426663 544070 426672
rect 543922 413264 543978 413273
rect 543922 413199 543978 413208
rect 543830 252104 543886 252113
rect 543830 252039 543886 252048
rect 543832 180600 543884 180606
rect 543830 180568 543832 180577
rect 543884 180568 543886 180577
rect 543830 180503 543886 180512
rect 543832 167272 543884 167278
rect 543830 167240 543832 167249
rect 543884 167240 543886 167249
rect 543830 167175 543886 167184
rect 543830 162480 543886 162489
rect 543830 162415 543886 162424
rect 543844 150521 543872 162415
rect 543830 150512 543886 150521
rect 543830 150447 543886 150456
rect 543830 139496 543886 139505
rect 543830 139431 543886 139440
rect 543844 131345 543872 139431
rect 543830 131336 543886 131345
rect 543830 131271 543886 131280
rect 543738 109032 543794 109041
rect 543738 108967 543794 108976
rect 543738 104272 543794 104281
rect 543738 104207 543794 104216
rect 543556 104168 543608 104174
rect 543556 104110 543608 104116
rect 543372 95192 543424 95198
rect 543372 95134 543424 95140
rect 543384 44198 543412 95134
rect 543462 86320 543518 86329
rect 543462 86255 543518 86264
rect 543372 44192 543424 44198
rect 543372 44134 543424 44140
rect 543280 42560 543332 42566
rect 543280 42502 543332 42508
rect 543476 42226 543504 86255
rect 543568 73234 543596 104110
rect 543752 95198 543780 104207
rect 543740 95192 543792 95198
rect 543740 95134 543792 95140
rect 543830 81968 543886 81977
rect 543830 81903 543886 81912
rect 543844 81462 543872 81903
rect 543832 81456 543884 81462
rect 543832 81398 543884 81404
rect 543738 77344 543794 77353
rect 543738 77279 543794 77288
rect 543648 75880 543700 75886
rect 543648 75822 543700 75828
rect 543556 73228 543608 73234
rect 543556 73170 543608 73176
rect 543660 44334 543688 75822
rect 543648 44328 543700 44334
rect 543648 44270 543700 44276
rect 543556 44192 543608 44198
rect 543556 44134 543608 44140
rect 543464 42220 543516 42226
rect 543464 42162 543516 42168
rect 543188 3732 543240 3738
rect 543188 3674 543240 3680
rect 543568 3602 543596 44134
rect 543752 42498 543780 77279
rect 543832 69012 543884 69018
rect 543832 68954 543884 68960
rect 543844 68513 543872 68954
rect 543830 68504 543886 68513
rect 543830 68439 543886 68448
rect 543832 64184 543884 64190
rect 543830 64152 543832 64161
rect 543884 64152 543886 64161
rect 543830 64087 543886 64096
rect 543832 59560 543884 59566
rect 543830 59528 543832 59537
rect 543884 59528 543886 59537
rect 543830 59463 543886 59472
rect 543830 55040 543886 55049
rect 543830 54975 543886 54984
rect 543844 53854 543872 54975
rect 543832 53848 543884 53854
rect 543832 53790 543884 53796
rect 543830 50688 543886 50697
rect 543830 50623 543886 50632
rect 543740 42492 543792 42498
rect 543740 42434 543792 42440
rect 543844 42294 543872 50623
rect 543936 44062 543964 413199
rect 544014 373008 544070 373017
rect 544014 372943 544070 372952
rect 543924 44056 543976 44062
rect 543924 43998 543976 44004
rect 543832 42288 543884 42294
rect 543832 42230 543884 42236
rect 544028 5506 544056 372943
rect 544120 369209 544148 628079
rect 544212 475969 544240 700266
rect 544844 691416 544896 691422
rect 544844 691358 544896 691364
rect 544290 661464 544346 661473
rect 544290 661399 544346 661408
rect 544304 655110 544332 661399
rect 544384 661360 544436 661366
rect 544384 661302 544436 661308
rect 544292 655104 544344 655110
rect 544292 655046 544344 655052
rect 544292 654968 544344 654974
rect 544292 654910 544344 654916
rect 544198 475960 544254 475969
rect 544198 475895 544254 475904
rect 544200 417784 544252 417790
rect 544198 417752 544200 417761
rect 544252 417752 544254 417761
rect 544198 417687 544254 417696
rect 544200 409080 544252 409086
rect 544200 409022 544252 409028
rect 544212 408785 544240 409022
rect 544198 408776 544254 408785
rect 544198 408711 544254 408720
rect 544198 381984 544254 381993
rect 544198 381919 544254 381928
rect 544106 369200 544162 369209
rect 544106 369135 544162 369144
rect 544106 368520 544162 368529
rect 544106 368455 544162 368464
rect 544016 5500 544068 5506
rect 544016 5442 544068 5448
rect 544120 5166 544148 368455
rect 544212 44130 544240 381919
rect 544304 323921 544332 654910
rect 544396 328273 544424 661302
rect 544568 661292 544620 661298
rect 544568 661234 544620 661240
rect 544476 659932 544528 659938
rect 544476 659874 544528 659880
rect 544488 332897 544516 659874
rect 544580 654974 544608 661234
rect 544752 661156 544804 661162
rect 544752 661098 544804 661104
rect 544660 659660 544712 659666
rect 544660 659602 544712 659608
rect 544672 659569 544700 659602
rect 544658 659560 544714 659569
rect 544658 659495 544714 659504
rect 544764 659410 544792 661098
rect 544672 659382 544792 659410
rect 544568 654968 544620 654974
rect 544568 654910 544620 654916
rect 544568 654832 544620 654838
rect 544568 654774 544620 654780
rect 544580 346225 544608 654774
rect 544672 547738 544700 659382
rect 544752 659320 544804 659326
rect 544752 659262 544804 659268
rect 544660 547732 544712 547738
rect 544660 547674 544712 547680
rect 544658 547632 544714 547641
rect 544658 547567 544714 547576
rect 544672 546514 544700 547567
rect 544660 546508 544712 546514
rect 544660 546450 544712 546456
rect 544660 535424 544712 535430
rect 544660 535366 544712 535372
rect 544672 534177 544700 535366
rect 544658 534168 544714 534177
rect 544658 534103 544714 534112
rect 544660 520872 544712 520878
rect 544658 520840 544660 520849
rect 544712 520840 544714 520849
rect 544658 520775 544714 520784
rect 544660 511896 544712 511902
rect 544658 511864 544660 511873
rect 544712 511864 544714 511873
rect 544658 511799 544714 511808
rect 544658 507376 544714 507385
rect 544658 507311 544714 507320
rect 544672 506530 544700 507311
rect 544660 506524 544712 506530
rect 544660 506466 544712 506472
rect 544660 493944 544712 493950
rect 544658 493912 544660 493921
rect 544712 493912 544714 493921
rect 544658 493847 544714 493856
rect 544660 489592 544712 489598
rect 544658 489560 544660 489569
rect 544712 489560 544714 489569
rect 544658 489495 544714 489504
rect 544658 466848 544714 466857
rect 544658 466783 544714 466792
rect 544672 466478 544700 466783
rect 544660 466472 544712 466478
rect 544660 466414 544712 466420
rect 544660 462664 544712 462670
rect 544658 462632 544660 462641
rect 544712 462632 544714 462641
rect 544658 462567 544714 462576
rect 544658 453520 544714 453529
rect 544658 453455 544714 453464
rect 544672 452674 544700 453455
rect 544660 452668 544712 452674
rect 544660 452610 544712 452616
rect 544660 449880 544712 449886
rect 544660 449822 544712 449828
rect 544672 449313 544700 449822
rect 544658 449304 544714 449313
rect 544658 449239 544714 449248
rect 544658 445768 544714 445777
rect 544658 445703 544714 445712
rect 544566 346216 544622 346225
rect 544566 346151 544622 346160
rect 544566 337104 544622 337113
rect 544566 337039 544622 337048
rect 544474 332888 544530 332897
rect 544474 332823 544530 332832
rect 544382 328264 544438 328273
rect 544382 328199 544438 328208
rect 544290 323912 544346 323921
rect 544290 323847 544346 323856
rect 544290 314800 544346 314809
rect 544290 314735 544346 314744
rect 544200 44124 544252 44130
rect 544200 44066 544252 44072
rect 544304 43450 544332 314735
rect 544382 310176 544438 310185
rect 544382 310111 544438 310120
rect 544292 43444 544344 43450
rect 544292 43386 544344 43392
rect 544396 42158 544424 310111
rect 544476 229832 544528 229838
rect 544474 229800 544476 229809
rect 544528 229800 544530 229809
rect 544474 229735 544530 229744
rect 544474 211712 544530 211721
rect 544474 211647 544530 211656
rect 544488 211206 544516 211647
rect 544476 211200 544528 211206
rect 544476 211142 544528 211148
rect 544474 191720 544530 191729
rect 544474 191655 544530 191664
rect 544488 189582 544516 191655
rect 544476 189576 544528 189582
rect 544476 189518 544528 189524
rect 544474 171456 544530 171465
rect 544474 171391 544530 171400
rect 544488 171290 544516 171391
rect 544476 171284 544528 171290
rect 544476 171226 544528 171232
rect 544474 122224 544530 122233
rect 544474 122159 544530 122168
rect 544488 44266 544516 122159
rect 544476 44260 544528 44266
rect 544476 44202 544528 44208
rect 544384 42152 544436 42158
rect 544384 42094 544436 42100
rect 544580 37942 544608 337039
rect 544672 149297 544700 445703
rect 544764 400330 544792 659262
rect 544856 646241 544884 691358
rect 545120 664488 545172 664494
rect 545120 664430 545172 664436
rect 544936 660340 544988 660346
rect 544936 660282 544988 660288
rect 544842 646232 544898 646241
rect 544842 646167 544898 646176
rect 544844 637560 544896 637566
rect 544844 637502 544896 637508
rect 544856 637265 544884 637502
rect 544842 637256 544898 637265
rect 544842 637191 544898 637200
rect 544844 630012 544896 630018
rect 544844 629954 544896 629960
rect 544856 623937 544884 629954
rect 544842 623928 544898 623937
rect 544842 623863 544898 623872
rect 544842 619168 544898 619177
rect 544842 619103 544898 619112
rect 544856 618322 544884 619103
rect 544844 618316 544896 618322
rect 544844 618258 544896 618264
rect 544844 606008 544896 606014
rect 544842 605976 544844 605985
rect 544896 605976 544898 605985
rect 544842 605911 544898 605920
rect 544842 601216 544898 601225
rect 544842 601151 544898 601160
rect 544856 400450 544884 601151
rect 544948 574818 544976 660282
rect 545028 660068 545080 660074
rect 545028 660010 545080 660016
rect 545040 574938 545068 660010
rect 545028 574932 545080 574938
rect 545028 574874 545080 574880
rect 544948 574790 545068 574818
rect 544936 574728 544988 574734
rect 544934 574696 544936 574705
rect 544988 574696 544990 574705
rect 544934 574631 544990 574640
rect 544936 574592 544988 574598
rect 544936 574534 544988 574540
rect 544948 570081 544976 574534
rect 544934 570072 544990 570081
rect 544934 570007 544990 570016
rect 544936 565820 544988 565826
rect 544936 565762 544988 565768
rect 544948 565729 544976 565762
rect 544934 565720 544990 565729
rect 544934 565655 544990 565664
rect 545040 561105 545068 574790
rect 545026 561096 545082 561105
rect 545026 561031 545082 561040
rect 544936 552152 544988 552158
rect 544934 552120 544936 552129
rect 544988 552120 544990 552129
rect 544934 552055 544990 552064
rect 544936 547732 544988 547738
rect 544936 547674 544988 547680
rect 544948 538801 544976 547674
rect 544934 538792 544990 538801
rect 544934 538727 544990 538736
rect 545026 516352 545082 516361
rect 545026 516287 545082 516296
rect 545040 516186 545068 516287
rect 545028 516180 545080 516186
rect 545028 516122 545080 516128
rect 545026 498400 545082 498409
rect 545026 498335 545082 498344
rect 545040 498234 545068 498335
rect 545028 498228 545080 498234
rect 545028 498170 545080 498176
rect 545028 485852 545080 485858
rect 545028 485794 545080 485800
rect 544936 440360 544988 440366
rect 544934 440328 544936 440337
rect 544988 440328 544990 440337
rect 544934 440263 544990 440272
rect 544936 405680 544988 405686
rect 544936 405622 544988 405628
rect 544948 404433 544976 405622
rect 544934 404424 544990 404433
rect 544934 404359 544990 404368
rect 544844 400444 544896 400450
rect 544844 400386 544896 400392
rect 544764 400302 544976 400330
rect 544844 400240 544896 400246
rect 544844 400182 544896 400188
rect 544752 400172 544804 400178
rect 544752 400114 544804 400120
rect 544764 400081 544792 400114
rect 544750 400072 544806 400081
rect 544750 400007 544806 400016
rect 544752 396024 544804 396030
rect 544752 395966 544804 395972
rect 544764 395457 544792 395966
rect 544750 395448 544806 395457
rect 544750 395383 544806 395392
rect 544750 390960 544806 390969
rect 544750 390895 544806 390904
rect 544764 390658 544792 390895
rect 544752 390652 544804 390658
rect 544752 390594 544804 390600
rect 544752 377528 544804 377534
rect 544750 377496 544752 377505
rect 544804 377496 544806 377505
rect 544750 377431 544806 377440
rect 544752 364200 544804 364206
rect 544750 364168 544752 364177
rect 544804 364168 544806 364177
rect 544750 364103 544806 364112
rect 544856 362982 544884 400182
rect 544948 397458 544976 400302
rect 544936 397452 544988 397458
rect 544936 397394 544988 397400
rect 545040 393314 545068 485794
rect 544948 393286 545068 393314
rect 544948 386481 544976 393286
rect 544934 386472 544990 386481
rect 544934 386407 544990 386416
rect 544844 362976 544896 362982
rect 544844 362918 544896 362924
rect 544934 359408 544990 359417
rect 544934 359343 544990 359352
rect 544948 358834 544976 359343
rect 544936 358828 544988 358834
rect 544936 358770 544988 358776
rect 544752 342236 544804 342242
rect 544752 342178 544804 342184
rect 544764 341873 544792 342178
rect 544750 341864 544806 341873
rect 544750 341799 544806 341808
rect 544934 319152 544990 319161
rect 544934 319087 544990 319096
rect 544948 318986 544976 319087
rect 544936 318980 544988 318986
rect 544936 318922 544988 318928
rect 544934 278896 544990 278905
rect 544934 278831 544990 278840
rect 544948 278798 544976 278831
rect 544936 278792 544988 278798
rect 544936 278734 544988 278740
rect 544752 275664 544804 275670
rect 544752 275606 544804 275612
rect 544764 274689 544792 275606
rect 544750 274680 544806 274689
rect 544750 274615 544806 274624
rect 544934 269920 544990 269929
rect 544934 269855 544990 269864
rect 544750 256592 544806 256601
rect 544750 256527 544806 256536
rect 544764 255338 544792 256527
rect 544752 255332 544804 255338
rect 544752 255274 544804 255280
rect 544750 247616 544806 247625
rect 544750 247551 544806 247560
rect 544764 247110 544792 247551
rect 544752 247104 544804 247110
rect 544752 247046 544804 247052
rect 544750 242992 544806 243001
rect 544750 242927 544752 242936
rect 544804 242927 544806 242936
rect 544752 242898 544804 242904
rect 544750 238640 544806 238649
rect 544750 238575 544806 238584
rect 544764 237454 544792 238575
rect 544752 237448 544804 237454
rect 544752 237390 544804 237396
rect 544750 225312 544806 225321
rect 544750 225247 544806 225256
rect 544764 225010 544792 225247
rect 544752 225004 544804 225010
rect 544752 224946 544804 224952
rect 544750 220688 544806 220697
rect 544750 220623 544806 220632
rect 544764 219502 544792 220623
rect 544752 219496 544804 219502
rect 544752 219438 544804 219444
rect 544752 208344 544804 208350
rect 544752 208286 544804 208292
rect 544764 207505 544792 208286
rect 544750 207496 544806 207505
rect 544750 207431 544806 207440
rect 544750 184784 544806 184793
rect 544750 184719 544806 184728
rect 544764 183598 544792 184719
rect 544752 183592 544804 183598
rect 544752 183534 544804 183540
rect 544752 176656 544804 176662
rect 544752 176598 544804 176604
rect 544764 175953 544792 176598
rect 544750 175944 544806 175953
rect 544750 175879 544806 175888
rect 544752 158704 544804 158710
rect 544752 158646 544804 158652
rect 544764 158273 544792 158646
rect 544750 158264 544806 158273
rect 544750 158199 544806 158208
rect 544658 149288 544714 149297
rect 544658 149223 544714 149232
rect 544660 114504 544712 114510
rect 544660 114446 544712 114452
rect 544672 113393 544700 114446
rect 544658 113384 544714 113393
rect 544658 113319 544714 113328
rect 544658 99920 544714 99929
rect 544658 99855 544714 99864
rect 544672 46986 544700 99855
rect 544750 90944 544806 90953
rect 544750 90879 544806 90888
rect 544660 46980 544712 46986
rect 544660 46922 544712 46928
rect 544660 46844 544712 46850
rect 544660 46786 544712 46792
rect 544672 46209 544700 46786
rect 544658 46200 544714 46209
rect 544658 46135 544714 46144
rect 544660 46096 544712 46102
rect 544660 46038 544712 46044
rect 544672 43382 544700 46038
rect 544764 44198 544792 90879
rect 544844 86284 544896 86290
rect 544844 86226 544896 86232
rect 544856 46102 544884 86226
rect 544844 46096 544896 46102
rect 544844 46038 544896 46044
rect 544844 45960 544896 45966
rect 544844 45902 544896 45908
rect 544752 44192 544804 44198
rect 544752 44134 544804 44140
rect 544856 43518 544884 45902
rect 544948 44402 544976 269855
rect 545026 126576 545082 126585
rect 545026 126511 545082 126520
rect 545040 45966 545068 126511
rect 545028 45960 545080 45966
rect 545028 45902 545080 45908
rect 545028 45824 545080 45830
rect 545028 45766 545080 45772
rect 544936 44396 544988 44402
rect 544936 44338 544988 44344
rect 544844 43512 544896 43518
rect 544844 43454 544896 43460
rect 544660 43376 544712 43382
rect 544660 43318 544712 43324
rect 545040 42362 545068 45766
rect 545028 42356 545080 42362
rect 545028 42298 545080 42304
rect 544568 37936 544620 37942
rect 544568 37878 544620 37884
rect 545132 6322 545160 664430
rect 545212 662040 545264 662046
rect 545212 661982 545264 661988
rect 545120 6316 545172 6322
rect 545120 6258 545172 6264
rect 544108 5160 544160 5166
rect 544108 5102 544160 5108
rect 543556 3596 543608 3602
rect 543556 3538 543608 3544
rect 543004 3324 543056 3330
rect 543004 3266 543056 3272
rect 545224 3262 545252 661982
rect 545316 660550 545344 702406
rect 547420 700460 547472 700466
rect 547420 700402 547472 700408
rect 546868 663740 546920 663746
rect 546868 663682 546920 663688
rect 546684 663468 546736 663474
rect 546684 663410 546736 663416
rect 545396 663332 545448 663338
rect 545396 663274 545448 663280
rect 545304 660544 545356 660550
rect 545304 660486 545356 660492
rect 545302 578368 545358 578377
rect 545302 578303 545358 578312
rect 545316 578270 545344 578303
rect 545304 578264 545356 578270
rect 545304 578206 545356 578212
rect 545302 556608 545358 556617
rect 545302 556543 545358 556552
rect 545316 42634 545344 556543
rect 545408 364206 545436 663274
rect 546500 663060 546552 663066
rect 546500 663002 546552 663008
rect 545672 662312 545724 662318
rect 545672 662254 545724 662260
rect 545488 662108 545540 662114
rect 545488 662050 545540 662056
rect 545500 431390 545528 662050
rect 545580 661768 545632 661774
rect 545580 661710 545632 661716
rect 545592 435742 545620 661710
rect 545684 489598 545712 662254
rect 545764 662176 545816 662182
rect 545764 662118 545816 662124
rect 545672 489592 545724 489598
rect 545672 489534 545724 489540
rect 545580 435736 545632 435742
rect 545580 435678 545632 435684
rect 545488 431384 545540 431390
rect 545488 431326 545540 431332
rect 545396 364200 545448 364206
rect 545396 364142 545448 364148
rect 545396 362976 545448 362982
rect 545396 362918 545448 362924
rect 545304 42628 545356 42634
rect 545304 42570 545356 42576
rect 545408 3534 545436 362918
rect 545670 287872 545726 287881
rect 545670 287807 545726 287816
rect 545486 265568 545542 265577
rect 545486 265503 545542 265512
rect 545500 5302 545528 265503
rect 545684 240106 545712 287807
rect 545672 240100 545724 240106
rect 545672 240042 545724 240048
rect 545578 216336 545634 216345
rect 545578 216271 545634 216280
rect 545488 5296 545540 5302
rect 545488 5238 545540 5244
rect 545592 5030 545620 216271
rect 545670 189408 545726 189417
rect 545670 189343 545726 189352
rect 545684 171834 545712 189343
rect 545672 171828 545724 171834
rect 545672 171770 545724 171776
rect 545776 81394 545804 662118
rect 545948 661904 546000 661910
rect 545948 661846 546000 661852
rect 545856 582412 545908 582418
rect 545856 582354 545908 582360
rect 545764 81388 545816 81394
rect 545764 81330 545816 81336
rect 545670 72992 545726 73001
rect 545670 72927 545726 72936
rect 545684 5438 545712 72927
rect 545868 40594 545896 582354
rect 545960 511902 545988 661846
rect 546040 547188 546092 547194
rect 546040 547130 546092 547136
rect 546052 537538 546080 547130
rect 546040 537532 546092 537538
rect 546040 537474 546092 537480
rect 546132 516180 546184 516186
rect 546132 516122 546184 516128
rect 545948 511896 546000 511902
rect 545948 511838 546000 511844
rect 545948 474768 546000 474774
rect 545948 474710 546000 474716
rect 545960 64190 545988 474710
rect 546040 380996 546092 381002
rect 546040 380938 546092 380944
rect 545948 64184 546000 64190
rect 545948 64126 546000 64132
rect 546052 43790 546080 380938
rect 546144 338094 546172 516122
rect 546132 338088 546184 338094
rect 546132 338030 546184 338036
rect 546408 336728 546460 336734
rect 546408 336670 546460 336676
rect 546132 316736 546184 316742
rect 546132 316678 546184 316684
rect 546144 43926 546172 316678
rect 546224 287700 546276 287706
rect 546224 287642 546276 287648
rect 546132 43920 546184 43926
rect 546132 43862 546184 43868
rect 546040 43784 546092 43790
rect 546040 43726 546092 43732
rect 546236 43178 546264 287642
rect 546316 267028 546368 267034
rect 546316 266970 546368 266976
rect 546328 43654 546356 266970
rect 546420 265742 546448 336670
rect 546408 265736 546460 265742
rect 546408 265678 546460 265684
rect 546408 189576 546460 189582
rect 546408 189518 546460 189524
rect 546420 184958 546448 189518
rect 546408 184952 546460 184958
rect 546408 184894 546460 184900
rect 546408 180872 546460 180878
rect 546408 180814 546460 180820
rect 546420 43858 546448 180814
rect 546512 59566 546540 663002
rect 546592 659728 546644 659734
rect 546592 659670 546644 659676
rect 546604 167278 546632 659670
rect 546696 180606 546724 663410
rect 546776 662380 546828 662386
rect 546776 662322 546828 662328
rect 546788 409086 546816 662322
rect 546880 417790 546908 663682
rect 547144 662788 547196 662794
rect 547144 662730 547196 662736
rect 546960 613420 547012 613426
rect 546960 613362 547012 613368
rect 546972 606014 547000 613362
rect 546960 606008 547012 606014
rect 546960 605950 547012 605956
rect 546868 417784 546920 417790
rect 546868 417726 546920 417732
rect 546776 409080 546828 409086
rect 546776 409022 546828 409028
rect 547050 291136 547106 291145
rect 547050 291071 547106 291080
rect 547064 265674 547092 291071
rect 547052 265668 547104 265674
rect 547052 265610 547104 265616
rect 546684 180600 546736 180606
rect 546684 180542 546736 180548
rect 546592 167272 546644 167278
rect 546592 167214 546644 167220
rect 546500 59560 546552 59566
rect 546500 59502 546552 59508
rect 546408 43852 546460 43858
rect 546408 43794 546460 43800
rect 546316 43648 546368 43654
rect 546316 43590 546368 43596
rect 546224 43172 546276 43178
rect 546224 43114 546276 43120
rect 545856 40588 545908 40594
rect 545856 40530 545908 40536
rect 547156 37262 547184 662730
rect 547328 661836 547380 661842
rect 547328 661778 547380 661784
rect 547236 572756 547288 572762
rect 547236 572698 547288 572704
rect 547248 41274 547276 572698
rect 547340 140758 547368 661778
rect 547432 229838 547460 700402
rect 547604 664760 547656 664766
rect 547604 664702 547656 664708
rect 547512 478916 547564 478922
rect 547512 478858 547564 478864
rect 547420 229832 547472 229838
rect 547420 229774 547472 229780
rect 547420 211200 547472 211206
rect 547420 211142 547472 211148
rect 547432 194546 547460 211142
rect 547420 194540 547472 194546
rect 547420 194482 547472 194488
rect 547420 171284 547472 171290
rect 547420 171226 547472 171232
rect 547328 140752 547380 140758
rect 547328 140694 547380 140700
rect 547236 41268 547288 41274
rect 547236 41210 547288 41216
rect 547144 37256 547196 37262
rect 547144 37198 547196 37204
rect 545672 5432 545724 5438
rect 545672 5374 545724 5380
rect 545580 5024 545632 5030
rect 545580 4966 545632 4972
rect 547432 4010 547460 171226
rect 547524 40458 547552 478858
rect 547616 460902 547644 664702
rect 547788 498228 547840 498234
rect 547788 498170 547840 498176
rect 547604 460896 547656 460902
rect 547604 460838 547656 460844
rect 547604 444440 547656 444446
rect 547604 444382 547656 444388
rect 547512 40452 547564 40458
rect 547512 40394 547564 40400
rect 547616 39778 547644 444382
rect 547696 331016 547748 331022
rect 547696 330958 547748 330964
rect 547708 322930 547736 330958
rect 547696 322924 547748 322930
rect 547696 322866 547748 322872
rect 547696 292596 547748 292602
rect 547696 292538 547748 292544
rect 547708 41410 547736 292538
rect 547800 284306 547828 498170
rect 547788 284300 547840 284306
rect 547788 284242 547840 284248
rect 547788 164280 547840 164286
rect 547788 164222 547840 164228
rect 547696 41404 547748 41410
rect 547696 41346 547748 41352
rect 547800 41342 547828 164222
rect 547788 41336 547840 41342
rect 547788 41278 547840 41284
rect 547604 39772 547656 39778
rect 547604 39714 547656 39720
rect 547892 38962 547920 703582
rect 548904 703474 548932 703582
rect 549046 703520 549158 704960
rect 552032 703582 552244 703610
rect 549088 703474 549116 703520
rect 548904 703446 549116 703474
rect 550180 700324 550232 700330
rect 550180 700266 550232 700272
rect 548524 666596 548576 666602
rect 548524 666538 548576 666544
rect 548340 386164 548392 386170
rect 548340 386106 548392 386112
rect 548352 381002 548380 386106
rect 548340 380996 548392 381002
rect 548340 380938 548392 380944
rect 548536 41138 548564 666538
rect 548892 664692 548944 664698
rect 548892 664634 548944 664640
rect 548708 664352 548760 664358
rect 548708 664294 548760 664300
rect 548616 662652 548668 662658
rect 548616 662594 548668 662600
rect 548628 180810 548656 662594
rect 548720 558890 548748 664294
rect 548800 664012 548852 664018
rect 548800 663954 548852 663960
rect 548708 558884 548760 558890
rect 548708 558826 548760 558832
rect 548708 538892 548760 538898
rect 548708 538834 548760 538840
rect 548720 520878 548748 538834
rect 548708 520872 548760 520878
rect 548708 520814 548760 520820
rect 548708 503736 548760 503742
rect 548708 503678 548760 503684
rect 548616 180804 548668 180810
rect 548616 180746 548668 180752
rect 548616 149116 548668 149122
rect 548616 149058 548668 149064
rect 548524 41132 548576 41138
rect 548524 41074 548576 41080
rect 548628 39098 548656 149058
rect 548616 39092 548668 39098
rect 548616 39034 548668 39040
rect 548720 39030 548748 503678
rect 548812 500954 548840 663954
rect 548904 579630 548932 664634
rect 549996 664420 550048 664426
rect 549996 664362 550048 664368
rect 549260 664148 549312 664154
rect 549260 664090 549312 664096
rect 548984 663944 549036 663950
rect 548984 663886 549036 663892
rect 548996 604450 549024 663886
rect 549076 660000 549128 660006
rect 549076 659942 549128 659948
rect 549088 623762 549116 659942
rect 549076 623756 549128 623762
rect 549076 623698 549128 623704
rect 548984 604444 549036 604450
rect 548984 604386 549036 604392
rect 548984 587920 549036 587926
rect 548984 587862 549036 587868
rect 548892 579624 548944 579630
rect 548892 579566 548944 579572
rect 548996 552158 549024 587862
rect 548984 552152 549036 552158
rect 548984 552094 549036 552100
rect 548800 500948 548852 500954
rect 548800 500890 548852 500896
rect 548800 484424 548852 484430
rect 548800 484366 548852 484372
rect 548812 462670 548840 484366
rect 548800 462664 548852 462670
rect 548800 462606 548852 462612
rect 548800 449948 548852 449954
rect 548800 449890 548852 449896
rect 548812 39846 548840 449890
rect 548892 425128 548944 425134
rect 548892 425070 548944 425076
rect 548904 40050 548932 425070
rect 548984 386436 549036 386442
rect 548984 386378 549036 386384
rect 548996 40934 549024 386378
rect 549076 196036 549128 196042
rect 549076 195978 549128 195984
rect 549088 180878 549116 195978
rect 549076 180872 549128 180878
rect 549076 180814 549128 180820
rect 549076 135312 549128 135318
rect 549076 135254 549128 135260
rect 548984 40928 549036 40934
rect 548984 40870 549036 40876
rect 548892 40044 548944 40050
rect 548892 39986 548944 39992
rect 548800 39840 548852 39846
rect 548800 39782 548852 39788
rect 549088 39642 549116 135254
rect 549076 39636 549128 39642
rect 549076 39578 549128 39584
rect 548708 39024 548760 39030
rect 548708 38966 548760 38972
rect 547880 38956 547932 38962
rect 547880 38898 547932 38904
rect 547420 4004 547472 4010
rect 547420 3946 547472 3952
rect 545396 3528 545448 3534
rect 545396 3470 545448 3476
rect 545212 3256 545264 3262
rect 545212 3198 545264 3204
rect 549272 480 549300 664090
rect 549904 616888 549956 616894
rect 549904 616830 549956 616836
rect 549352 501628 549404 501634
rect 549352 501570 549404 501576
rect 549364 493950 549392 501570
rect 549352 493944 549404 493950
rect 549352 493886 549404 493892
rect 549812 184884 549864 184890
rect 549812 184826 549864 184832
rect 549824 178090 549852 184826
rect 549812 178084 549864 178090
rect 549812 178026 549864 178032
rect 549536 79824 549588 79830
rect 549536 79766 549588 79772
rect 549548 75954 549576 79766
rect 549536 75948 549588 75954
rect 549536 75890 549588 75896
rect 549916 39302 549944 616830
rect 550008 102134 550036 664362
rect 550088 641776 550140 641782
rect 550088 641718 550140 641724
rect 550100 597038 550128 641718
rect 550088 597032 550140 597038
rect 550088 596974 550140 596980
rect 550088 454096 550140 454102
rect 550088 454038 550140 454044
rect 550100 440366 550128 454038
rect 550088 440360 550140 440366
rect 550088 440302 550140 440308
rect 550088 434784 550140 434790
rect 550088 434726 550140 434732
rect 549996 102128 550048 102134
rect 549996 102070 550048 102076
rect 550100 39506 550128 434726
rect 550192 377534 550220 700266
rect 552032 665854 552060 703582
rect 552216 703474 552244 703582
rect 552358 703520 552470 704960
rect 555670 703520 555782 704960
rect 558982 703520 559094 704960
rect 562294 703520 562406 704960
rect 564452 703582 565492 703610
rect 552400 703474 552428 703520
rect 552216 703446 552428 703474
rect 555712 700466 555740 703520
rect 555700 700460 555752 700466
rect 555700 700402 555752 700408
rect 552756 685908 552808 685914
rect 552756 685850 552808 685856
rect 552020 665848 552072 665854
rect 552020 665790 552072 665796
rect 551284 665100 551336 665106
rect 551284 665042 551336 665048
rect 550272 663876 550324 663882
rect 550272 663818 550324 663824
rect 550180 377528 550232 377534
rect 550180 377470 550232 377476
rect 550284 376718 550312 663818
rect 550364 607232 550416 607238
rect 550364 607174 550416 607180
rect 550376 574734 550404 607174
rect 550364 574728 550416 574734
rect 550364 574670 550416 574676
rect 550456 528624 550508 528630
rect 550456 528566 550508 528572
rect 550364 397452 550416 397458
rect 550364 397394 550416 397400
rect 550376 391270 550404 397394
rect 550364 391264 550416 391270
rect 550364 391206 550416 391212
rect 550272 376712 550324 376718
rect 550272 376654 550324 376660
rect 550180 356108 550232 356114
rect 550180 356050 550232 356056
rect 550088 39500 550140 39506
rect 550088 39442 550140 39448
rect 549904 39296 549956 39302
rect 549904 39238 549956 39244
rect 550192 38826 550220 356050
rect 550272 318980 550324 318986
rect 550272 318922 550324 318928
rect 550284 307766 550312 318922
rect 550272 307760 550324 307766
rect 550272 307702 550324 307708
rect 550272 302252 550324 302258
rect 550272 302194 550324 302200
rect 550180 38820 550232 38826
rect 550180 38762 550232 38768
rect 550284 38758 550312 302194
rect 550364 296744 550416 296750
rect 550364 296686 550416 296692
rect 550376 39574 550404 296686
rect 550468 275670 550496 528566
rect 550824 488572 550876 488578
rect 550824 488514 550876 488520
rect 550836 482225 550864 488514
rect 550822 482216 550878 482225
rect 550822 482151 550878 482160
rect 551192 390856 551244 390862
rect 551192 390798 551244 390804
rect 551204 386170 551232 390798
rect 551192 386164 551244 386170
rect 551192 386106 551244 386112
rect 550548 382628 550600 382634
rect 550548 382570 550600 382576
rect 550560 378146 550588 382570
rect 550548 378140 550600 378146
rect 550548 378082 550600 378088
rect 550548 287088 550600 287094
rect 550548 287030 550600 287036
rect 550456 275664 550508 275670
rect 550456 275606 550508 275612
rect 550456 255332 550508 255338
rect 550456 255274 550508 255280
rect 550468 175234 550496 255274
rect 550456 175228 550508 175234
rect 550456 175170 550508 175176
rect 550364 39568 550416 39574
rect 550364 39510 550416 39516
rect 550560 38894 550588 287030
rect 551192 237448 551244 237454
rect 551192 237390 551244 237396
rect 551100 205692 551152 205698
rect 551100 205634 551152 205640
rect 551112 196042 551140 205634
rect 551100 196036 551152 196042
rect 551100 195978 551152 195984
rect 551204 131102 551232 237390
rect 551192 131096 551244 131102
rect 551192 131038 551244 131044
rect 551192 84244 551244 84250
rect 551192 84186 551244 84192
rect 551204 79830 551232 84186
rect 551192 79824 551244 79830
rect 551192 79766 551244 79772
rect 550548 38888 550600 38894
rect 550548 38830 550600 38836
rect 550272 38752 550324 38758
rect 550272 38694 550324 38700
rect 551296 3534 551324 665042
rect 551376 664624 551428 664630
rect 551376 664566 551428 664572
rect 551388 27606 551416 664566
rect 551836 664284 551888 664290
rect 551836 664226 551888 664232
rect 551560 664216 551612 664222
rect 551560 664158 551612 664164
rect 551468 661156 551520 661162
rect 551468 661098 551520 661104
rect 551480 39914 551508 661098
rect 551572 46918 551600 664158
rect 551652 494080 551704 494086
rect 551652 494022 551704 494028
rect 551560 46912 551612 46918
rect 551560 46854 551612 46860
rect 551468 39908 551520 39914
rect 551468 39850 551520 39856
rect 551664 39681 551692 494022
rect 551744 440292 551796 440298
rect 551744 440234 551796 440240
rect 551756 396030 551784 440234
rect 551744 396024 551796 396030
rect 551744 395966 551796 395972
rect 551744 390584 551796 390590
rect 551744 390526 551796 390532
rect 551650 39672 551706 39681
rect 551650 39607 551706 39616
rect 551756 39438 551784 390526
rect 551848 372570 551876 664226
rect 552662 664048 552718 664057
rect 552662 663983 552718 663992
rect 552572 409896 552624 409902
rect 552572 409838 552624 409844
rect 552584 405686 552612 409838
rect 552572 405680 552624 405686
rect 552572 405622 552624 405628
rect 551928 390652 551980 390658
rect 551928 390594 551980 390600
rect 551836 372564 551888 372570
rect 551836 372506 551888 372512
rect 551836 365764 551888 365770
rect 551836 365706 551888 365712
rect 551744 39432 551796 39438
rect 551744 39374 551796 39380
rect 551848 39166 551876 365706
rect 551940 313274 551968 390594
rect 552572 378140 552624 378146
rect 552572 378082 552624 378088
rect 552584 374950 552612 378082
rect 552572 374944 552624 374950
rect 552572 374886 552624 374892
rect 551928 313268 551980 313274
rect 551928 313210 551980 313216
rect 551928 258120 551980 258126
rect 551928 258062 551980 258068
rect 551940 39710 551968 258062
rect 552020 45552 552072 45558
rect 552020 45494 552072 45500
rect 552032 44169 552060 45494
rect 552018 44160 552074 44169
rect 552018 44095 552074 44104
rect 551928 39704 551980 39710
rect 551928 39646 551980 39652
rect 551836 39160 551888 39166
rect 551836 39102 551888 39108
rect 551376 27600 551428 27606
rect 551376 27542 551428 27548
rect 552676 3534 552704 663983
rect 552768 41206 552796 685850
rect 559024 683114 559052 703520
rect 562336 700330 562364 703520
rect 562324 700324 562376 700330
rect 562324 700266 562376 700272
rect 558932 683086 559052 683114
rect 554044 670744 554096 670750
rect 554044 670686 554096 670692
rect 553032 664896 553084 664902
rect 553032 664838 553084 664844
rect 552848 664080 552900 664086
rect 552848 664022 552900 664028
rect 552860 184890 552888 664022
rect 552940 469260 552992 469266
rect 552940 469202 552992 469208
rect 552848 184884 552900 184890
rect 552848 184826 552900 184832
rect 552848 120148 552900 120154
rect 552848 120090 552900 120096
rect 552756 41200 552808 41206
rect 552756 41142 552808 41148
rect 552860 38690 552888 120090
rect 552952 39982 552980 469202
rect 553044 278730 553072 664838
rect 553400 537532 553452 537538
rect 553400 537474 553452 537480
rect 553412 533390 553440 537474
rect 554056 535430 554084 670686
rect 558932 664562 558960 683086
rect 558920 664556 558972 664562
rect 558920 664498 558972 664504
rect 562322 653440 562378 653449
rect 562322 653375 562378 653384
rect 562336 651438 562364 653375
rect 562324 651432 562376 651438
rect 562324 651374 562376 651380
rect 563704 636268 563756 636274
rect 563704 636210 563756 636216
rect 558276 600976 558328 600982
rect 558276 600918 558328 600924
rect 558184 597576 558236 597582
rect 558184 597518 558236 597524
rect 556804 553444 556856 553450
rect 556804 553386 556856 553392
rect 554044 535424 554096 535430
rect 554044 535366 554096 535372
rect 553400 533384 553452 533390
rect 553400 533326 553452 533332
rect 554136 506524 554188 506530
rect 554136 506466 554188 506472
rect 554044 489932 554096 489938
rect 554044 489874 554096 489880
rect 553124 405748 553176 405754
rect 553124 405690 553176 405696
rect 553136 400178 553164 405690
rect 553124 400172 553176 400178
rect 553124 400114 553176 400120
rect 553308 346452 553360 346458
rect 553308 346394 553360 346400
rect 553320 342242 553348 346394
rect 553308 342236 553360 342242
rect 553308 342178 553360 342184
rect 553124 299600 553176 299606
rect 553124 299542 553176 299548
rect 553136 287706 553164 299542
rect 553124 287700 553176 287706
rect 553124 287642 553176 287648
rect 553308 278792 553360 278798
rect 553308 278734 553360 278740
rect 553032 278724 553084 278730
rect 553032 278666 553084 278672
rect 553320 274650 553348 278734
rect 553308 274644 553360 274650
rect 553308 274586 553360 274592
rect 553032 270768 553084 270774
rect 553032 270710 553084 270716
rect 553044 267034 553072 270710
rect 553032 267028 553084 267034
rect 553032 266970 553084 266976
rect 553032 247104 553084 247110
rect 553032 247046 553084 247052
rect 553044 234598 553072 247046
rect 553032 234592 553084 234598
rect 553032 234534 553084 234540
rect 553124 225004 553176 225010
rect 553124 224946 553176 224952
rect 553032 219496 553084 219502
rect 553032 219438 553084 219444
rect 553044 200122 553072 219438
rect 553136 209778 553164 224946
rect 553124 209772 553176 209778
rect 553124 209714 553176 209720
rect 553400 209092 553452 209098
rect 553400 209034 553452 209040
rect 553412 205698 553440 209034
rect 553400 205692 553452 205698
rect 553400 205634 553452 205640
rect 553032 200116 553084 200122
rect 553032 200058 553084 200064
rect 554056 69018 554084 489874
rect 554148 190466 554176 506466
rect 556160 302388 556212 302394
rect 556160 302330 556212 302336
rect 556172 299606 556200 302330
rect 556160 299600 556212 299606
rect 556160 299542 556212 299548
rect 554780 273964 554832 273970
rect 554780 273906 554832 273912
rect 554792 270774 554820 273906
rect 554780 270768 554832 270774
rect 554780 270710 554832 270716
rect 554136 190460 554188 190466
rect 554136 190402 554188 190408
rect 554688 178016 554740 178022
rect 554688 177958 554740 177964
rect 554700 175250 554728 177958
rect 554700 175222 554820 175250
rect 554792 172990 554820 175222
rect 554780 172984 554832 172990
rect 554780 172926 554832 172932
rect 556816 158710 556844 553386
rect 557540 395344 557592 395350
rect 557540 395286 557592 395292
rect 557552 390862 557580 395286
rect 557540 390856 557592 390862
rect 557540 390798 557592 390804
rect 556896 265736 556948 265742
rect 556896 265678 556948 265684
rect 556908 251870 556936 265678
rect 556896 251864 556948 251870
rect 556896 251806 556948 251812
rect 556804 158704 556856 158710
rect 556804 158646 556856 158652
rect 558196 114510 558224 597518
rect 558288 597514 558316 600918
rect 558276 597508 558328 597514
rect 558276 597450 558328 597456
rect 562968 597508 563020 597514
rect 562968 597450 563020 597456
rect 562980 593366 563008 597450
rect 562968 593360 563020 593366
rect 562968 593302 563020 593308
rect 562324 546508 562376 546514
rect 562324 546450 562376 546456
rect 559564 538280 559616 538286
rect 559564 538222 559616 538228
rect 558920 492380 558972 492386
rect 558920 492322 558972 492328
rect 558932 488578 558960 492322
rect 558920 488572 558972 488578
rect 558920 488514 558972 488520
rect 558368 374944 558420 374950
rect 558368 374886 558420 374892
rect 558276 352572 558328 352578
rect 558276 352514 558328 352520
rect 558288 316742 558316 352514
rect 558380 350198 558408 374886
rect 558368 350192 558420 350198
rect 558368 350134 558420 350140
rect 558276 316736 558328 316742
rect 558276 316678 558328 316684
rect 559576 176662 559604 538222
rect 561036 466472 561088 466478
rect 561036 466414 561088 466420
rect 560944 358828 560996 358834
rect 560944 358770 560996 358776
rect 559656 311160 559708 311166
rect 559656 311102 559708 311108
rect 559668 302394 559696 311102
rect 559656 302388 559708 302394
rect 559656 302330 559708 302336
rect 560956 219434 560984 358770
rect 561048 353258 561076 466414
rect 562048 458856 562100 458862
rect 562048 458798 562100 458804
rect 562060 455462 562088 458798
rect 562048 455456 562100 455462
rect 562048 455398 562100 455404
rect 562336 401606 562364 546450
rect 562324 401600 562376 401606
rect 562324 401542 562376 401548
rect 563060 391264 563112 391270
rect 563060 391206 563112 391212
rect 563072 388482 563100 391206
rect 563060 388476 563112 388482
rect 563060 388418 563112 388424
rect 561036 353252 561088 353258
rect 561036 353194 561088 353200
rect 561036 350192 561088 350198
rect 561036 350134 561088 350140
rect 561048 340882 561076 350134
rect 561036 340876 561088 340882
rect 561036 340818 561088 340824
rect 563336 287700 563388 287706
rect 563336 287642 563388 287648
rect 563348 284374 563376 287642
rect 561036 284368 561088 284374
rect 561036 284310 561088 284316
rect 563336 284368 563388 284374
rect 563336 284310 563388 284316
rect 561048 273970 561076 284310
rect 561036 273964 561088 273970
rect 561036 273906 561088 273912
rect 563060 265668 563112 265674
rect 563060 265610 563112 265616
rect 563072 260166 563100 265610
rect 563060 260160 563112 260166
rect 563060 260102 563112 260108
rect 561036 242956 561088 242962
rect 561036 242898 561088 242904
rect 560944 219428 560996 219434
rect 560944 219370 560996 219376
rect 559564 176656 559616 176662
rect 559564 176598 559616 176604
rect 558920 172984 558972 172990
rect 558920 172926 558972 172932
rect 558932 170406 558960 172926
rect 558920 170400 558972 170406
rect 558920 170342 558972 170348
rect 561048 117298 561076 242898
rect 561036 117292 561088 117298
rect 561036 117234 561088 117240
rect 558184 114504 558236 114510
rect 558184 114446 558236 114452
rect 561772 89752 561824 89758
rect 561772 89694 561824 89700
rect 561784 85610 561812 89694
rect 558828 85604 558880 85610
rect 558828 85546 558880 85552
rect 561772 85604 561824 85610
rect 561772 85546 561824 85552
rect 558840 84250 558868 85546
rect 558828 84244 558880 84250
rect 558828 84186 558880 84192
rect 558184 81456 558236 81462
rect 558184 81398 558236 81404
rect 554044 69012 554096 69018
rect 554044 68954 554096 68960
rect 554778 43616 554834 43625
rect 554778 43551 554834 43560
rect 552940 39976 552992 39982
rect 552940 39918 552992 39924
rect 552848 38684 552900 38690
rect 552848 38626 552900 38632
rect 554792 16574 554820 43551
rect 558196 42770 558224 81398
rect 559840 47524 559892 47530
rect 559840 47466 559892 47472
rect 559852 45626 559880 47466
rect 563716 46850 563744 636210
rect 563796 507136 563848 507142
rect 563796 507078 563848 507084
rect 563808 492386 563836 507078
rect 563796 492380 563848 492386
rect 563796 492322 563848 492328
rect 564452 208350 564480 703582
rect 565464 703474 565492 703582
rect 565606 703520 565718 704960
rect 568592 703582 568804 703610
rect 565648 703474 565676 703520
rect 565464 703446 565676 703474
rect 565820 661088 565872 661094
rect 565820 661030 565872 661036
rect 565084 533384 565136 533390
rect 565084 533326 565136 533332
rect 565096 527134 565124 533326
rect 565084 527128 565136 527134
rect 565084 527070 565136 527076
rect 564440 208344 564492 208350
rect 564440 208286 564492 208292
rect 565084 183592 565136 183598
rect 565084 183534 565136 183540
rect 565096 155922 565124 183534
rect 565084 155916 565136 155922
rect 565084 155858 565136 155864
rect 563796 94512 563848 94518
rect 563796 94454 563848 94460
rect 563808 86290 563836 94454
rect 563796 86284 563848 86290
rect 563796 86226 563848 86232
rect 564440 52828 564492 52834
rect 564440 52770 564492 52776
rect 564452 47530 564480 52770
rect 564440 47524 564492 47530
rect 564440 47466 564492 47472
rect 563704 46844 563756 46850
rect 563704 46786 563756 46792
rect 559840 45620 559892 45626
rect 559840 45562 559892 45568
rect 558184 42764 558236 42770
rect 558184 42706 558236 42712
rect 554792 16546 555464 16574
rect 551284 3528 551336 3534
rect 551284 3470 551336 3476
rect 552572 3528 552624 3534
rect 552572 3470 552624 3476
rect 552664 3528 552716 3534
rect 552664 3470 552716 3476
rect 552584 480 552612 3470
rect 555436 490 555464 16546
rect 559196 3800 559248 3806
rect 559196 3742 559248 3748
rect 555712 598 555924 626
rect 555712 490 555740 598
rect 539110 -960 539222 480
rect 542422 -960 542534 480
rect 545734 -960 545846 480
rect 549230 -960 549342 480
rect 552542 -960 552654 480
rect 555436 462 555740 490
rect 555896 480 555924 598
rect 559208 480 559236 3742
rect 562508 3392 562560 3398
rect 562508 3334 562560 3340
rect 562520 480 562548 3334
rect 565832 480 565860 661030
rect 568592 660482 568620 703582
rect 568776 703474 568804 703582
rect 568918 703520 569030 704960
rect 571352 703582 572116 703610
rect 568960 703474 568988 703520
rect 568776 703446 568988 703474
rect 568580 660476 568632 660482
rect 568580 660418 568632 660424
rect 567844 651364 567896 651370
rect 567844 651306 567896 651312
rect 567856 648650 567884 651306
rect 567844 648644 567896 648650
rect 567844 648586 567896 648592
rect 567844 578264 567896 578270
rect 567844 578206 567896 578212
rect 566464 455456 566516 455462
rect 566464 455398 566516 455404
rect 566476 442270 566504 455398
rect 566464 442264 566516 442270
rect 566464 442206 566516 442212
rect 567752 110492 567804 110498
rect 567752 110434 567804 110440
rect 567764 104174 567792 110434
rect 567752 104168 567804 104174
rect 567752 104110 567804 104116
rect 566464 97300 566516 97306
rect 566464 97242 566516 97248
rect 566476 89758 566504 97242
rect 566464 89752 566516 89758
rect 566464 89694 566516 89700
rect 567856 52426 567884 578206
rect 569040 527128 569092 527134
rect 569040 527070 569092 527076
rect 569052 522986 569080 527070
rect 569040 522980 569092 522986
rect 569040 522922 569092 522928
rect 569868 398132 569920 398138
rect 569868 398074 569920 398080
rect 569880 395350 569908 398074
rect 569868 395344 569920 395350
rect 569868 395286 569920 395292
rect 570604 388476 570656 388482
rect 570604 388418 570656 388424
rect 570616 382226 570644 388418
rect 570604 382220 570656 382226
rect 570604 382162 570656 382168
rect 569224 340876 569276 340882
rect 569224 340818 569276 340824
rect 569236 334422 569264 340818
rect 569224 334416 569276 334422
rect 569224 334358 569276 334364
rect 570604 223304 570656 223310
rect 570604 223246 570656 223252
rect 570616 209098 570644 223246
rect 570604 209092 570656 209098
rect 570604 209034 570656 209040
rect 569684 170400 569736 170406
rect 569684 170342 569736 170348
rect 569696 167074 569724 170342
rect 569684 167068 569736 167074
rect 569684 167010 569736 167016
rect 567936 59356 567988 59362
rect 567936 59298 567988 59304
rect 567948 52834 567976 59298
rect 567936 52828 567988 52834
rect 567936 52770 567988 52776
rect 567844 52420 567896 52426
rect 567844 52362 567896 52368
rect 571352 41002 571380 703582
rect 572088 703474 572116 703582
rect 572230 703520 572342 704960
rect 575542 703520 575654 704960
rect 578854 703520 578966 704960
rect 581012 703582 582052 703610
rect 572272 703474 572300 703520
rect 572088 703446 572300 703474
rect 575584 701010 575612 703520
rect 575572 701004 575624 701010
rect 575572 700946 575624 700952
rect 578896 700398 578924 703520
rect 578884 700392 578936 700398
rect 578884 700334 578936 700340
rect 580630 696416 580686 696425
rect 580630 696351 580686 696360
rect 580170 691520 580226 691529
rect 580170 691455 580226 691464
rect 580184 691422 580212 691455
rect 580172 691416 580224 691422
rect 580172 691358 580224 691364
rect 579618 686624 579674 686633
rect 579618 686559 579674 686568
rect 579632 685914 579660 686559
rect 579620 685908 579672 685914
rect 579620 685850 579672 685856
rect 580170 681728 580226 681737
rect 580170 681663 580226 681672
rect 580184 680406 580212 681663
rect 580172 680400 580224 680406
rect 580172 680342 580224 680348
rect 580170 671936 580226 671945
rect 580170 671871 580226 671880
rect 580184 670750 580212 671871
rect 580172 670744 580224 670750
rect 580172 670686 580224 670692
rect 579618 667040 579674 667049
rect 579618 666975 579674 666984
rect 579632 666602 579660 666975
rect 579620 666596 579672 666602
rect 579620 666538 579672 666544
rect 580448 663604 580500 663610
rect 580448 663546 580500 663552
rect 580356 662720 580408 662726
rect 580356 662662 580408 662668
rect 579618 662144 579674 662153
rect 579618 662079 579674 662088
rect 579632 661162 579660 662079
rect 580264 661972 580316 661978
rect 580264 661914 580316 661920
rect 579620 661156 579672 661162
rect 579620 661098 579672 661104
rect 580172 659796 580224 659802
rect 580172 659738 580224 659744
rect 571984 648576 572036 648582
rect 571984 648518 572036 648524
rect 571996 629270 572024 648518
rect 580078 642288 580134 642297
rect 580078 642223 580134 642232
rect 580092 641782 580120 642223
rect 580080 641776 580132 641782
rect 580080 641718 580132 641724
rect 579986 637392 580042 637401
rect 579986 637327 580042 637336
rect 580000 636274 580028 637327
rect 579988 636268 580040 636274
rect 579988 636210 580040 636216
rect 580184 632505 580212 659738
rect 580170 632496 580226 632505
rect 580170 632431 580226 632440
rect 571984 629264 572036 629270
rect 571984 629206 572036 629212
rect 575480 629264 575532 629270
rect 575480 629206 575532 629212
rect 575492 626618 575520 629206
rect 575480 626612 575532 626618
rect 575480 626554 575532 626560
rect 576860 626612 576912 626618
rect 576860 626554 576912 626560
rect 576872 621518 576900 626554
rect 580172 623756 580224 623762
rect 580172 623698 580224 623704
rect 580184 622713 580212 623698
rect 580170 622704 580226 622713
rect 580170 622639 580226 622648
rect 576860 621512 576912 621518
rect 576860 621454 576912 621460
rect 579528 621512 579580 621518
rect 579528 621454 579580 621460
rect 578884 618316 578936 618322
rect 578884 618258 578936 618264
rect 571984 522980 572036 522986
rect 571984 522922 572036 522928
rect 571996 518226 572024 522922
rect 577504 521212 577556 521218
rect 577504 521154 577556 521160
rect 571984 518220 572036 518226
rect 571984 518162 572036 518168
rect 577516 509318 577544 521154
rect 574100 509312 574152 509318
rect 574100 509254 574152 509260
rect 577504 509312 577556 509318
rect 577504 509254 577556 509260
rect 574112 507142 574140 509254
rect 574100 507136 574152 507142
rect 574100 507078 574152 507084
rect 574744 452668 574796 452674
rect 574744 452610 574796 452616
rect 574100 442264 574152 442270
rect 574100 442206 574152 442212
rect 574112 437442 574140 442206
rect 574100 437436 574152 437442
rect 574100 437378 574152 437384
rect 574100 334416 574152 334422
rect 574100 334358 574152 334364
rect 574112 328438 574140 334358
rect 574100 328432 574152 328438
rect 574100 328374 574152 328380
rect 572720 251864 572772 251870
rect 572720 251806 572772 251812
rect 572732 249762 572760 251806
rect 572720 249756 572772 249762
rect 572720 249698 572772 249704
rect 574008 229152 574060 229158
rect 574008 229094 574060 229100
rect 574020 223310 574048 229094
rect 574008 223304 574060 223310
rect 574008 223246 574060 223252
rect 574756 215286 574784 452610
rect 577504 437436 577556 437442
rect 577504 437378 577556 437384
rect 577516 431458 577544 437378
rect 577504 431452 577556 431458
rect 577504 431394 577556 431400
rect 574836 361616 574888 361622
rect 574836 361558 574888 361564
rect 574848 352578 574876 361558
rect 574836 352572 574888 352578
rect 574836 352514 574888 352520
rect 575480 313948 575532 313954
rect 575480 313890 575532 313896
rect 575492 311166 575520 313890
rect 575480 311160 575532 311166
rect 575480 311102 575532 311108
rect 577504 302320 577556 302326
rect 577504 302262 577556 302268
rect 577516 287706 577544 302262
rect 577504 287700 577556 287706
rect 577504 287642 577556 287648
rect 574744 215280 574796 215286
rect 574744 215222 574796 215228
rect 574744 167000 574796 167006
rect 574744 166942 574796 166948
rect 574756 160138 574784 166942
rect 574744 160132 574796 160138
rect 574744 160074 574796 160080
rect 578240 102196 578292 102202
rect 578240 102138 578292 102144
rect 578252 100858 578280 102138
rect 578160 100830 578280 100858
rect 578160 97306 578188 100830
rect 578148 97300 578200 97306
rect 578148 97242 578200 97248
rect 578896 86329 578924 618258
rect 579540 618202 579568 621454
rect 579540 618174 579660 618202
rect 579632 612921 579660 618174
rect 579986 617808 580042 617817
rect 579986 617743 580042 617752
rect 580000 616894 580028 617743
rect 579988 616888 580040 616894
rect 579988 616830 580040 616836
rect 579618 612912 579674 612921
rect 579618 612847 579674 612856
rect 580170 608016 580226 608025
rect 580170 607951 580226 607960
rect 580184 607238 580212 607951
rect 580172 607232 580224 607238
rect 580172 607174 580224 607180
rect 579620 604444 579672 604450
rect 579620 604386 579672 604392
rect 579632 603129 579660 604386
rect 579618 603120 579674 603129
rect 579618 603055 579674 603064
rect 580170 598224 580226 598233
rect 580170 598159 580226 598168
rect 580184 597582 580212 598159
rect 580172 597576 580224 597582
rect 580172 597518 580224 597524
rect 579620 593360 579672 593366
rect 579620 593302 579672 593308
rect 579632 593065 579660 593302
rect 579618 593056 579674 593065
rect 579618 592991 579674 593000
rect 580170 588160 580226 588169
rect 580170 588095 580226 588104
rect 580184 587926 580212 588095
rect 580172 587920 580224 587926
rect 580172 587862 580224 587868
rect 579986 583264 580042 583273
rect 579986 583199 580042 583208
rect 580000 582418 580028 583199
rect 579988 582412 580040 582418
rect 579988 582354 580040 582360
rect 579620 579624 579672 579630
rect 579620 579566 579672 579572
rect 579632 578377 579660 579566
rect 579618 578368 579674 578377
rect 579618 578303 579674 578312
rect 580170 573472 580226 573481
rect 580170 573407 580226 573416
rect 580184 572762 580212 573407
rect 580172 572756 580224 572762
rect 580172 572698 580224 572704
rect 580172 558884 580224 558890
rect 580172 558826 580224 558832
rect 580184 558793 580212 558826
rect 580170 558784 580226 558793
rect 580170 558719 580226 558728
rect 580170 553888 580226 553897
rect 580170 553823 580226 553832
rect 580184 553450 580212 553823
rect 580172 553444 580224 553450
rect 580172 553386 580224 553392
rect 580078 544096 580134 544105
rect 580078 544031 580134 544040
rect 580092 538898 580120 544031
rect 580170 538928 580226 538937
rect 580080 538892 580132 538898
rect 580170 538863 580226 538872
rect 580080 538834 580132 538840
rect 580184 538286 580212 538863
rect 580172 538280 580224 538286
rect 580172 538222 580224 538228
rect 580276 534041 580304 661914
rect 580262 534032 580318 534041
rect 580262 533967 580318 533976
rect 580170 529136 580226 529145
rect 580170 529071 580226 529080
rect 580184 528630 580212 529071
rect 580172 528624 580224 528630
rect 580172 528566 580224 528572
rect 579618 524240 579674 524249
rect 579618 524175 579674 524184
rect 579632 521218 579660 524175
rect 579620 521212 579672 521218
rect 579620 521154 579672 521160
rect 580262 519344 580318 519353
rect 580262 519279 580318 519288
rect 580172 518220 580224 518226
rect 580172 518162 580224 518168
rect 580184 514457 580212 518162
rect 580170 514448 580226 514457
rect 580170 514383 580226 514392
rect 579986 504656 580042 504665
rect 579986 504591 580042 504600
rect 580000 503742 580028 504591
rect 579988 503736 580040 503742
rect 579988 503678 580040 503684
rect 579712 500948 579764 500954
rect 579712 500890 579764 500896
rect 579724 499769 579752 500890
rect 579710 499760 579766 499769
rect 579710 499695 579766 499704
rect 579986 494864 580042 494873
rect 579986 494799 580042 494808
rect 580000 494086 580028 494799
rect 579988 494080 580040 494086
rect 579988 494022 580040 494028
rect 580170 489968 580226 489977
rect 580170 489903 580172 489912
rect 580224 489903 580226 489912
rect 580172 489874 580224 489880
rect 580170 484800 580226 484809
rect 580170 484735 580226 484744
rect 580184 484430 580212 484735
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579618 479904 579674 479913
rect 579618 479839 579674 479848
rect 579632 478922 579660 479839
rect 579620 478916 579672 478922
rect 579620 478858 579672 478864
rect 580170 475008 580226 475017
rect 580170 474943 580226 474952
rect 580184 474774 580212 474943
rect 580172 474768 580224 474774
rect 580172 474710 580224 474716
rect 579986 470112 580042 470121
rect 579986 470047 580042 470056
rect 580000 469266 580028 470047
rect 579988 469260 580040 469266
rect 579988 469202 580040 469208
rect 580172 460896 580224 460902
rect 580172 460838 580224 460844
rect 580184 460329 580212 460838
rect 580170 460320 580226 460329
rect 580170 460255 580226 460264
rect 580170 455424 580226 455433
rect 580170 455359 580226 455368
rect 580184 454102 580212 455359
rect 580172 454096 580224 454102
rect 580172 454038 580224 454044
rect 580170 450528 580226 450537
rect 580170 450463 580226 450472
rect 580184 449954 580212 450463
rect 580172 449948 580224 449954
rect 580172 449890 580224 449896
rect 580170 445632 580226 445641
rect 580170 445567 580226 445576
rect 580184 444446 580212 445567
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 580170 440736 580226 440745
rect 580170 440671 580226 440680
rect 580184 440298 580212 440671
rect 580172 440292 580224 440298
rect 580172 440234 580224 440240
rect 580170 435840 580226 435849
rect 580170 435775 580226 435784
rect 580184 434790 580212 435775
rect 580172 434784 580224 434790
rect 580172 434726 580224 434732
rect 579620 431452 579672 431458
rect 579620 431394 579672 431400
rect 579632 430681 579660 431394
rect 579618 430672 579674 430681
rect 579618 430607 579674 430616
rect 580170 425776 580226 425785
rect 580170 425711 580226 425720
rect 580184 425134 580212 425711
rect 580172 425128 580224 425134
rect 580172 425070 580224 425076
rect 580170 411088 580226 411097
rect 580170 411023 580226 411032
rect 580184 409902 580212 411023
rect 580172 409896 580224 409902
rect 580172 409838 580224 409844
rect 580170 406192 580226 406201
rect 580170 406127 580226 406136
rect 580184 405754 580212 406127
rect 580172 405748 580224 405754
rect 580172 405690 580224 405696
rect 579712 401600 579764 401606
rect 579712 401542 579764 401548
rect 579724 401305 579752 401542
rect 579710 401296 579766 401305
rect 579710 401231 579766 401240
rect 579618 391504 579674 391513
rect 579618 391439 579674 391448
rect 579632 390590 579660 391439
rect 579620 390584 579672 390590
rect 579620 390526 579672 390532
rect 580170 386608 580226 386617
rect 580170 386543 580226 386552
rect 580184 386442 580212 386543
rect 580172 386436 580224 386442
rect 580172 386378 580224 386384
rect 579804 382220 579856 382226
rect 579804 382162 579856 382168
rect 579816 381721 579844 382162
rect 579802 381712 579858 381721
rect 579802 381647 579858 381656
rect 580172 376712 580224 376718
rect 580172 376654 580224 376660
rect 580184 376553 580212 376654
rect 580170 376544 580226 376553
rect 580170 376479 580226 376488
rect 579620 372564 579672 372570
rect 579620 372506 579672 372512
rect 579632 371657 579660 372506
rect 579618 371648 579674 371657
rect 579618 371583 579674 371592
rect 580170 366752 580226 366761
rect 580170 366687 580226 366696
rect 580184 365770 580212 366687
rect 580172 365764 580224 365770
rect 580172 365706 580224 365712
rect 580170 361856 580226 361865
rect 580170 361791 580226 361800
rect 580184 361622 580212 361791
rect 580172 361616 580224 361622
rect 580172 361558 580224 361564
rect 579986 356960 580042 356969
rect 579986 356895 580042 356904
rect 580000 356114 580028 356895
rect 579988 356108 580040 356114
rect 579988 356050 580040 356056
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 352073 580212 353194
rect 580170 352064 580226 352073
rect 580170 351999 580226 352008
rect 580170 347168 580226 347177
rect 580170 347103 580226 347112
rect 580184 346458 580212 347103
rect 580172 346452 580224 346458
rect 580172 346394 580224 346400
rect 580172 338088 580224 338094
rect 580172 338030 580224 338036
rect 580184 337385 580212 338030
rect 580170 337376 580226 337385
rect 580170 337311 580226 337320
rect 579988 328432 580040 328438
rect 579988 328374 580040 328380
rect 580000 327593 580028 328374
rect 579986 327584 580042 327593
rect 579986 327519 580042 327528
rect 579804 322924 579856 322930
rect 579804 322866 579856 322872
rect 579816 322425 579844 322866
rect 579802 322416 579858 322425
rect 579802 322351 579858 322360
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312633 580212 313210
rect 580170 312624 580226 312633
rect 580170 312559 580226 312568
rect 580172 307760 580224 307766
rect 580170 307728 580172 307737
rect 580224 307728 580226 307737
rect 580170 307663 580226 307672
rect 580170 302832 580226 302841
rect 580170 302767 580226 302776
rect 580184 302258 580212 302767
rect 580172 302252 580224 302258
rect 580172 302194 580224 302200
rect 579618 297936 579674 297945
rect 579618 297871 579674 297880
rect 579632 296750 579660 297871
rect 579620 296744 579672 296750
rect 579620 296686 579672 296692
rect 579802 293040 579858 293049
rect 579802 292975 579858 292984
rect 579816 292602 579844 292975
rect 579804 292596 579856 292602
rect 579804 292538 579856 292544
rect 579618 288144 579674 288153
rect 579618 288079 579674 288088
rect 579632 287094 579660 288079
rect 579620 287088 579672 287094
rect 579620 287030 579672 287036
rect 579620 284300 579672 284306
rect 579620 284242 579672 284248
rect 579632 283257 579660 284242
rect 579618 283248 579674 283257
rect 579618 283183 579674 283192
rect 579988 278724 580040 278730
rect 579988 278666 580040 278672
rect 580000 278361 580028 278666
rect 579986 278352 580042 278361
rect 579986 278287 580042 278296
rect 580172 274644 580224 274650
rect 580172 274586 580224 274592
rect 580184 273465 580212 274586
rect 580170 273456 580226 273465
rect 580170 273391 580226 273400
rect 579804 260160 579856 260166
rect 579804 260102 579856 260108
rect 579816 253609 579844 260102
rect 580170 258496 580226 258505
rect 580170 258431 580226 258440
rect 580184 258126 580212 258431
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 579802 253600 579858 253609
rect 579802 253535 579858 253544
rect 579620 249756 579672 249762
rect 579620 249698 579672 249704
rect 579632 248713 579660 249698
rect 579618 248704 579674 248713
rect 579618 248639 579674 248648
rect 580172 240100 580224 240106
rect 580172 240042 580224 240048
rect 580184 238921 580212 240042
rect 580170 238912 580226 238921
rect 580170 238847 580226 238856
rect 579988 234592 580040 234598
rect 579988 234534 580040 234540
rect 580000 234025 580028 234534
rect 579986 234016 580042 234025
rect 579986 233951 580042 233960
rect 580172 229152 580224 229158
rect 580170 229120 580172 229129
rect 580224 229120 580226 229129
rect 580170 229055 580226 229064
rect 579804 219428 579856 219434
rect 579804 219370 579856 219376
rect 579816 219337 579844 219370
rect 579802 219328 579858 219337
rect 579802 219263 579858 219272
rect 580172 215280 580224 215286
rect 580172 215222 580224 215228
rect 580184 214169 580212 215222
rect 580170 214160 580226 214169
rect 580170 214095 580226 214104
rect 579988 209772 580040 209778
rect 579988 209714 580040 209720
rect 580000 209273 580028 209714
rect 579986 209264 580042 209273
rect 579986 209199 580042 209208
rect 580172 200116 580224 200122
rect 580172 200058 580224 200064
rect 580184 199481 580212 200058
rect 580170 199472 580226 199481
rect 580170 199407 580226 199416
rect 580170 194576 580226 194585
rect 580170 194511 580172 194520
rect 580224 194511 580226 194520
rect 580172 194482 580224 194488
rect 579620 190460 579672 190466
rect 579620 190402 579672 190408
rect 579632 189689 579660 190402
rect 579618 189680 579674 189689
rect 579618 189615 579674 189624
rect 580172 184884 580224 184890
rect 580172 184826 580224 184832
rect 580184 184793 580212 184826
rect 580170 184784 580226 184793
rect 580170 184719 580226 184728
rect 579988 180804 580040 180810
rect 579988 180746 580040 180752
rect 580000 179897 580028 180746
rect 579986 179888 580042 179897
rect 579986 179823 580042 179832
rect 579620 175228 579672 175234
rect 579620 175170 579672 175176
rect 579632 175001 579660 175170
rect 579618 174992 579674 175001
rect 579618 174927 579674 174936
rect 579986 165200 580042 165209
rect 579986 165135 580042 165144
rect 580000 164286 580028 165135
rect 579988 164280 580040 164286
rect 579988 164222 580040 164228
rect 580172 160064 580224 160070
rect 580170 160032 580172 160041
rect 580224 160032 580226 160041
rect 580170 159967 580226 159976
rect 579620 155916 579672 155922
rect 579620 155858 579672 155864
rect 579632 155145 579660 155858
rect 579618 155136 579674 155145
rect 579618 155071 579674 155080
rect 579618 150240 579674 150249
rect 579618 150175 579674 150184
rect 579632 149122 579660 150175
rect 579620 149116 579672 149122
rect 579620 149058 579672 149064
rect 580172 140752 580224 140758
rect 580172 140694 580224 140700
rect 580184 140457 580212 140694
rect 580170 140448 580226 140457
rect 580170 140383 580226 140392
rect 579618 135552 579674 135561
rect 579618 135487 579674 135496
rect 579632 135318 579660 135487
rect 579620 135312 579672 135318
rect 579620 135254 579672 135260
rect 579804 131096 579856 131102
rect 579804 131038 579856 131044
rect 579816 130665 579844 131038
rect 579802 130656 579858 130665
rect 579802 130591 579858 130600
rect 580170 120864 580226 120873
rect 580170 120799 580226 120808
rect 580184 120154 580212 120799
rect 580172 120148 580224 120154
rect 580172 120090 580224 120096
rect 579620 117292 579672 117298
rect 579620 117234 579672 117240
rect 579632 115977 579660 117234
rect 579618 115968 579674 115977
rect 579618 115903 579674 115912
rect 580170 111072 580226 111081
rect 580170 111007 580226 111016
rect 580184 110498 580212 111007
rect 580172 110492 580224 110498
rect 580172 110434 580224 110440
rect 580170 105904 580226 105913
rect 580170 105839 580226 105848
rect 580184 102202 580212 105839
rect 580172 102196 580224 102202
rect 580172 102138 580224 102144
rect 579620 102128 579672 102134
rect 579620 102070 579672 102076
rect 579632 101017 579660 102070
rect 579618 101008 579674 101017
rect 579618 100943 579674 100952
rect 578974 96112 579030 96121
rect 578974 96047 579030 96056
rect 578882 86320 578938 86329
rect 578882 86255 578938 86264
rect 578988 66298 579016 96047
rect 580170 81424 580226 81433
rect 580170 81359 580172 81368
rect 580224 81359 580226 81368
rect 580172 81330 580224 81336
rect 575480 66292 575532 66298
rect 575480 66234 575532 66240
rect 578976 66292 579028 66298
rect 578976 66234 579028 66240
rect 575492 64874 575520 66234
rect 575400 64846 575520 64874
rect 575400 62150 575428 64846
rect 575388 62144 575440 62150
rect 575388 62086 575440 62092
rect 571708 62076 571760 62082
rect 571708 62018 571760 62024
rect 571720 59362 571748 62018
rect 580170 61840 580226 61849
rect 580170 61775 580226 61784
rect 571708 59356 571760 59362
rect 571708 59298 571760 59304
rect 580078 56944 580134 56953
rect 580078 56879 580134 56888
rect 579988 52420 580040 52426
rect 579988 52362 580040 52368
rect 580000 51785 580028 52362
rect 579986 51776 580042 51785
rect 579986 51711 580042 51720
rect 579988 46912 580040 46918
rect 579986 46880 579988 46889
rect 580040 46880 580042 46889
rect 579986 46815 580042 46824
rect 580092 44538 580120 56879
rect 580080 44532 580132 44538
rect 580080 44474 580132 44480
rect 580184 42922 580212 61775
rect 580092 42894 580212 42922
rect 571340 40996 571392 41002
rect 571340 40938 571392 40944
rect 580092 40390 580120 42894
rect 580172 42764 580224 42770
rect 580172 42706 580224 42712
rect 580184 41993 580212 42706
rect 580170 41984 580226 41993
rect 580170 41919 580226 41928
rect 580080 40384 580132 40390
rect 580080 40326 580132 40332
rect 580276 39370 580304 519279
rect 580368 243817 580396 662662
rect 580460 268297 580488 663546
rect 580540 661564 580592 661570
rect 580540 661506 580592 661512
rect 580552 549001 580580 661506
rect 580644 660414 580672 696351
rect 580906 676832 580962 676841
rect 580906 676767 580962 676776
rect 580724 661700 580776 661706
rect 580724 661642 580776 661648
rect 580632 660408 580684 660414
rect 580632 660350 580684 660356
rect 580630 652352 580686 652361
rect 580630 652287 580686 652296
rect 580644 565826 580672 652287
rect 580632 565820 580684 565826
rect 580632 565762 580684 565768
rect 580538 548992 580594 549001
rect 580538 548927 580594 548936
rect 580538 509552 580594 509561
rect 580538 509487 580594 509496
rect 580552 501634 580580 509487
rect 580540 501628 580592 501634
rect 580540 501570 580592 501576
rect 580538 465216 580594 465225
rect 580538 465151 580594 465160
rect 580552 449886 580580 465151
rect 580540 449880 580592 449886
rect 580540 449822 580592 449828
rect 580630 420880 580686 420889
rect 580630 420815 580686 420824
rect 580538 415984 580594 415993
rect 580538 415919 580594 415928
rect 580446 268288 580502 268297
rect 580446 268223 580502 268232
rect 580446 263392 580502 263401
rect 580446 263327 580502 263336
rect 580354 243808 580410 243817
rect 580354 243743 580410 243752
rect 580354 204368 580410 204377
rect 580354 204303 580410 204312
rect 580368 41070 580396 204303
rect 580460 44470 580488 263327
rect 580552 45554 580580 415919
rect 580644 398138 580672 420815
rect 580632 398132 580684 398138
rect 580632 398074 580684 398080
rect 580630 396400 580686 396409
rect 580630 396335 580686 396344
rect 580644 55214 580672 396335
rect 580736 342281 580764 661642
rect 580814 657248 580870 657257
rect 580814 657183 580870 657192
rect 580828 613426 580856 657183
rect 580920 637566 580948 676767
rect 581012 659666 581040 703582
rect 582024 703474 582052 703582
rect 582166 703520 582278 704960
rect 582208 703474 582236 703520
rect 582024 703446 582236 703474
rect 581000 659660 581052 659666
rect 581000 659602 581052 659608
rect 580908 637560 580960 637566
rect 580908 637502 580960 637508
rect 580816 613420 580868 613426
rect 580816 613362 580868 613368
rect 580722 342272 580778 342281
rect 580722 342207 580778 342216
rect 580722 332480 580778 332489
rect 580722 332415 580778 332424
rect 580736 313954 580764 332415
rect 580814 317520 580870 317529
rect 580814 317455 580870 317464
rect 580724 313948 580776 313954
rect 580724 313890 580776 313896
rect 580828 302326 580856 317455
rect 580816 302320 580868 302326
rect 580816 302262 580868 302268
rect 580908 171828 580960 171834
rect 580908 171770 580960 171776
rect 580920 170105 580948 171770
rect 580906 170096 580962 170105
rect 580906 170031 580962 170040
rect 580722 125760 580778 125769
rect 580722 125695 580778 125704
rect 580736 94518 580764 125695
rect 580724 94512 580776 94518
rect 580724 94454 580776 94460
rect 580814 71632 580870 71641
rect 580814 71567 580870 71576
rect 580644 55186 580764 55214
rect 580552 45526 580672 45554
rect 580540 44804 580592 44810
rect 580540 44746 580592 44752
rect 580448 44464 580500 44470
rect 580448 44406 580500 44412
rect 580448 42084 580500 42090
rect 580448 42026 580500 42032
rect 580356 41064 580408 41070
rect 580356 41006 580408 41012
rect 580264 39364 580316 39370
rect 580264 39306 580316 39312
rect 580172 37256 580224 37262
rect 580172 37198 580224 37204
rect 580184 37097 580212 37198
rect 580170 37088 580226 37097
rect 580170 37023 580226 37032
rect 580080 33108 580132 33114
rect 580080 33050 580132 33056
rect 580092 32201 580120 33050
rect 580078 32192 580134 32201
rect 580078 32127 580134 32136
rect 580080 27600 580132 27606
rect 580080 27542 580132 27548
rect 580092 27305 580120 27542
rect 580078 27296 580134 27305
rect 580078 27231 580134 27240
rect 580460 22409 580488 42026
rect 580552 40322 580580 44746
rect 580644 40526 580672 45526
rect 580736 44810 580764 55186
rect 580724 44804 580776 44810
rect 580724 44746 580776 44752
rect 580722 44704 580778 44713
rect 580722 44639 580778 44648
rect 580632 40520 580684 40526
rect 580632 40462 580684 40468
rect 580540 40316 580592 40322
rect 580540 40258 580592 40264
rect 580446 22400 580502 22409
rect 580446 22335 580502 22344
rect 580736 12617 580764 44639
rect 580828 40662 580856 71567
rect 580906 66736 580962 66745
rect 580906 66671 580962 66680
rect 580920 44606 580948 66671
rect 580908 44600 580960 44606
rect 580908 44542 580960 44548
rect 580816 40656 580868 40662
rect 580816 40598 580868 40604
rect 580722 12608 580778 12617
rect 580722 12543 580778 12552
rect 580172 8288 580224 8294
rect 580172 8230 580224 8236
rect 580184 7721 580212 8230
rect 580170 7712 580226 7721
rect 580170 7647 580226 7656
rect 575756 4140 575808 4146
rect 575756 4082 575808 4088
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 572444 3460 572496 3466
rect 572444 3402 572496 3408
rect 572456 480 572484 3402
rect 575768 480 575796 4082
rect 579068 4072 579120 4078
rect 579068 4014 579120 4020
rect 579080 480 579108 4014
rect 580172 4004 580224 4010
rect 580172 3946 580224 3952
rect 580184 2825 580212 3946
rect 582380 3868 582432 3874
rect 582380 3810 582432 3816
rect 580170 2816 580226 2825
rect 580170 2751 580226 2760
rect 582392 480 582420 3810
rect 555854 -960 555966 480
rect 559166 -960 559278 480
rect 562478 -960 562590 480
rect 565790 -960 565902 480
rect 569102 -960 569214 480
rect 572414 -960 572526 480
rect 575726 -960 575838 480
rect 579038 -960 579150 480
rect 582350 -960 582462 480
<< via2 >>
rect 3422 703704 3478 703760
rect 3238 698536 3294 698592
rect 3146 693640 3202 693696
rect 3514 688744 3570 688800
rect 3422 683848 3478 683904
rect 3422 664264 3478 664320
rect 3422 659368 3478 659424
rect 3422 654492 3478 654528
rect 3422 654472 3424 654492
rect 3424 654472 3476 654492
rect 3476 654472 3478 654492
rect 3330 649576 3386 649632
rect 2778 639512 2834 639568
rect 2778 634616 2834 634672
rect 3330 615032 3386 615088
rect 3330 610156 3386 610192
rect 3330 610136 3332 610156
rect 3332 610136 3384 610156
rect 3384 610136 3386 610156
rect 3330 605240 3386 605296
rect 2778 600344 2834 600400
rect 3330 595448 3386 595504
rect 3146 590316 3148 590336
rect 3148 590316 3200 590336
rect 3200 590316 3202 590336
rect 3146 590280 3202 590316
rect 2778 585384 2834 585440
rect 3238 580488 3294 580544
rect 3146 575592 3202 575648
rect 3054 570696 3110 570752
rect 2778 565800 2834 565856
rect 3146 560904 3202 560960
rect 3146 556008 3202 556064
rect 3146 551112 3202 551168
rect 3146 546216 3202 546272
rect 3146 541320 3202 541376
rect 2778 531276 2834 531312
rect 2778 531256 2780 531276
rect 2780 531256 2832 531276
rect 2832 531256 2834 531276
rect 3146 521464 3202 521520
rect 3146 511672 3202 511728
rect 3146 487192 3202 487248
rect 3054 482024 3110 482080
rect 2962 477128 3018 477184
rect 3146 467356 3202 467392
rect 3146 467336 3148 467356
rect 3148 467336 3200 467356
rect 3200 467336 3202 467356
rect 3146 462460 3202 462496
rect 3146 462440 3148 462460
rect 3148 462440 3200 462460
rect 3200 462440 3202 462460
rect 3238 457544 3294 457600
rect 3238 452648 3294 452704
rect 3146 447752 3202 447808
rect 3238 442856 3294 442912
rect 3238 437960 3294 438016
rect 2962 433064 3018 433120
rect 3238 427896 3294 427952
rect 3238 423000 3294 423056
rect 3238 418124 3294 418160
rect 3238 418104 3240 418124
rect 3240 418104 3292 418124
rect 3292 418104 3294 418124
rect 3146 413208 3202 413264
rect 2778 408348 2780 408368
rect 2780 408348 2832 408368
rect 2832 408348 2834 408368
rect 2778 408312 2834 408348
rect 3238 403416 3294 403472
rect 3238 398556 3240 398576
rect 3240 398556 3292 398576
rect 3292 398556 3294 398576
rect 3238 398520 3294 398556
rect 2778 393644 2834 393680
rect 2778 393624 2780 393644
rect 2780 393624 2832 393644
rect 2832 393624 2834 393644
rect 2778 383832 2834 383888
rect 3238 368872 3294 368928
rect 3330 363976 3386 364032
rect 3146 354184 3202 354240
rect 2778 349288 2834 349344
rect 3330 344412 3386 344448
rect 3330 344392 3332 344412
rect 3332 344392 3384 344412
rect 3384 344392 3386 344412
rect 3330 339516 3386 339552
rect 3330 339496 3332 339516
rect 3332 339496 3384 339516
rect 3384 339496 3386 339516
rect 2962 334600 3018 334656
rect 3238 329704 3294 329760
rect 3330 319640 3386 319696
rect 3330 314744 3386 314800
rect 2962 309848 3018 309904
rect 2778 304988 2780 305008
rect 2780 304988 2832 305008
rect 2832 304988 2834 305008
rect 2778 304952 2834 304988
rect 3330 300056 3386 300112
rect 3330 295160 3386 295216
rect 3146 290264 3202 290320
rect 3238 285368 3294 285424
rect 3146 265512 3202 265568
rect 3146 260616 3202 260672
rect 3146 226364 3202 226400
rect 3146 226344 3148 226364
rect 3148 226344 3200 226364
rect 3200 226344 3202 226364
rect 3054 216552 3110 216608
rect 3146 201592 3202 201648
rect 3146 196716 3202 196752
rect 3146 196696 3148 196716
rect 3148 196696 3200 196716
rect 3200 196696 3202 196716
rect 3146 186904 3202 186960
rect 3146 182008 3202 182064
rect 3054 177112 3110 177168
rect 3054 172216 3110 172272
rect 3146 167320 3202 167376
rect 2778 162460 2780 162480
rect 2780 162460 2832 162480
rect 2832 162460 2834 162480
rect 2778 162424 2834 162460
rect 2778 142568 2834 142624
rect 3330 280492 3386 280528
rect 3330 280472 3332 280492
rect 3332 280472 3384 280492
rect 3384 280472 3386 280492
rect 3330 275576 3386 275632
rect 3330 270680 3386 270736
rect 3238 127880 3294 127936
rect 3054 113212 3110 113248
rect 3054 113192 3056 113212
rect 3056 113192 3108 113212
rect 3108 113192 3110 113212
rect 3882 678952 3938 679008
rect 3698 674056 3754 674112
rect 3514 629720 3570 629776
rect 3790 669160 3846 669216
rect 3698 644408 3754 644464
rect 3882 624824 3938 624880
rect 3698 516568 3754 516624
rect 3514 506776 3570 506832
rect 3514 492088 3570 492144
rect 3514 472232 3570 472288
rect 3422 157256 3478 157312
rect 3422 147464 3478 147520
rect 3422 137672 3478 137728
rect 3422 132776 3478 132832
rect 3146 108296 3202 108352
rect 3330 103128 3386 103184
rect 2778 93336 2834 93392
rect 3330 83544 3386 83600
rect 2778 78684 2780 78704
rect 2780 78684 2832 78704
rect 2832 78684 2834 78704
rect 2778 78648 2834 78684
rect 3330 73752 3386 73808
rect 3330 68892 3332 68912
rect 3332 68892 3384 68912
rect 3384 68892 3386 68912
rect 3330 68856 3386 68892
rect 2778 63996 2780 64016
rect 2780 63996 2832 64016
rect 2832 63996 2834 64016
rect 2778 63960 2834 63996
rect 3330 54168 3386 54224
rect 2778 49000 2834 49056
rect 2778 39208 2834 39264
rect 3698 501880 3754 501936
rect 3698 496984 3754 497040
rect 3606 255720 3662 255776
rect 3606 245928 3662 245984
rect 3606 241068 3608 241088
rect 3608 241068 3660 241088
rect 3660 241068 3662 241088
rect 3606 241032 3662 241068
rect 3606 236172 3608 236192
rect 3608 236172 3660 236192
rect 3660 236172 3662 236192
rect 3606 236136 3662 236172
rect 3606 211384 3662 211440
rect 3790 250824 3846 250880
rect 3974 388728 4030 388784
rect 3974 373768 4030 373824
rect 3882 231240 3938 231296
rect 3882 221448 3938 221504
rect 3790 206488 3846 206544
rect 3882 191800 3938 191856
rect 3606 123004 3662 123040
rect 3606 122984 3608 123004
rect 3608 122984 3660 123004
rect 3660 122984 3662 123004
rect 3606 118088 3662 118144
rect 3606 88440 3662 88496
rect 3238 38936 3294 38992
rect 3422 34348 3424 34368
rect 3424 34348 3476 34368
rect 3476 34348 3478 34368
rect 3422 34312 3478 34348
rect 3238 24520 3294 24576
rect 3790 59064 3846 59120
rect 4066 359080 4122 359136
rect 4066 324808 4122 324864
rect 3882 43424 3938 43480
rect 4066 44104 4122 44160
rect 3882 29416 3938 29472
rect 3698 19624 3754 19680
rect 3422 14728 3478 14784
rect 2962 9868 2964 9888
rect 2964 9868 3016 9888
rect 3016 9868 3018 9888
rect 2962 9832 3018 9868
rect 6274 661136 6330 661192
rect 6182 40296 6238 40352
rect 8942 664808 8998 664864
rect 10322 40160 10378 40216
rect 10966 660184 11022 660240
rect 10506 40024 10562 40080
rect 10966 44512 11022 44568
rect 2778 4936 2834 4992
rect 35162 660728 35218 660784
rect 23386 39616 23442 39672
rect 38014 543360 38070 543416
rect 38014 520920 38070 520976
rect 37922 480664 37978 480720
rect 38106 122576 38162 122632
rect 38198 68720 38254 68776
rect 38106 44376 38162 44432
rect 38750 659776 38806 659832
rect 38658 565664 38714 565720
rect 38658 561312 38714 561368
rect 38658 556824 38714 556880
rect 38658 539008 38714 539064
rect 38658 529932 38660 529952
rect 38660 529932 38712 529952
rect 38712 529932 38714 529952
rect 38658 529896 38714 529932
rect 38658 525408 38714 525464
rect 38658 512080 38714 512136
rect 38842 655424 38898 655480
rect 38842 650800 38898 650856
rect 38842 646448 38898 646504
rect 38842 641824 38898 641880
rect 38934 628360 38990 628416
rect 38842 619384 38898 619440
rect 38842 615032 38898 615088
rect 38842 601604 38844 601624
rect 38844 601604 38896 601624
rect 38896 601604 38898 601624
rect 38842 601568 38898 601604
rect 38842 597216 38898 597272
rect 38842 592456 38898 592512
rect 38842 588240 38898 588296
rect 39026 579264 39082 579320
rect 38842 574504 38898 574560
rect 39118 570288 39174 570344
rect 38750 503104 38806 503160
rect 38750 498752 38806 498808
rect 38750 494128 38806 494184
rect 38750 489640 38806 489696
rect 38750 485152 38806 485208
rect 39394 660592 39450 660648
rect 39302 657328 39358 657384
rect 39210 547984 39266 548040
rect 39118 471824 39174 471880
rect 39302 467200 39358 467256
rect 38750 462848 38806 462904
rect 38750 458224 38806 458280
rect 38750 444760 38806 444816
rect 39302 435920 39358 435976
rect 38750 431568 38806 431624
rect 38750 426808 38806 426864
rect 39486 453872 39542 453928
rect 39394 422592 39450 422648
rect 38750 413480 38806 413536
rect 38750 399880 38806 399936
rect 39394 377712 39450 377768
rect 39394 373224 39450 373280
rect 38750 350648 38806 350704
rect 38750 346452 38806 346488
rect 38750 346432 38752 346452
rect 38752 346432 38804 346452
rect 38804 346432 38806 346452
rect 38750 332696 38806 332752
rect 38750 324128 38806 324184
rect 39302 319368 39358 319424
rect 38750 315016 38806 315072
rect 38750 310548 38806 310584
rect 38750 310528 38752 310548
rect 38752 310528 38804 310548
rect 38804 310528 38806 310548
rect 38750 306176 38806 306232
rect 38750 292576 38806 292632
rect 38750 283600 38806 283656
rect 39302 279248 39358 279304
rect 38750 270272 38806 270328
rect 38750 252184 38806 252240
rect 38842 247968 38898 248024
rect 38750 243344 38806 243400
rect 38750 238992 38806 239048
rect 38750 234368 38806 234424
rect 38750 229880 38806 229936
rect 38842 220904 38898 220960
rect 38842 207712 38898 207768
rect 39762 637472 39818 637528
rect 39762 582392 39818 582448
rect 39670 395664 39726 395720
rect 39578 391040 39634 391096
rect 39578 368600 39634 368656
rect 39670 341672 39726 341728
rect 39578 288088 39634 288144
rect 39486 203088 39542 203144
rect 38842 193976 38898 194032
rect 39486 189760 39542 189816
rect 38842 185000 38898 185056
rect 39118 180784 39174 180840
rect 38842 176160 38898 176216
rect 38842 167184 38898 167240
rect 38842 162696 38898 162752
rect 38934 140392 38990 140448
rect 38842 131552 38898 131608
rect 38842 113600 38898 113656
rect 38842 108996 38898 109032
rect 38842 108976 38844 108996
rect 38844 108976 38896 108996
rect 38896 108976 38898 108996
rect 39486 171672 39542 171728
rect 39302 158072 39358 158128
rect 39210 144744 39266 144800
rect 39026 95512 39082 95568
rect 38934 91160 38990 91216
rect 38842 86536 38898 86592
rect 38842 59608 38898 59664
rect 38842 43968 38898 44024
rect 39118 82184 39174 82240
rect 39394 135768 39450 135824
rect 39762 265920 39818 265976
rect 39946 632848 40002 632904
rect 39946 552336 40002 552392
rect 39946 534384 40002 534440
rect 39946 449248 40002 449304
rect 39854 261296 39910 261352
rect 39762 198736 39818 198792
rect 39946 153720 40002 153776
rect 40130 583616 40186 583672
rect 40130 507320 40186 507376
rect 40038 149504 40094 149560
rect 40038 126792 40094 126848
rect 39854 104488 39910 104544
rect 39946 99864 40002 99920
rect 40038 77560 40094 77616
rect 39854 73208 39910 73264
rect 39946 64232 40002 64288
rect 40222 440408 40278 440464
rect 40406 301552 40462 301608
rect 40406 297064 40462 297120
rect 40314 225392 40370 225448
rect 40314 216280 40370 216336
rect 40958 660456 41014 660512
rect 40590 328480 40646 328536
rect 40498 274624 40554 274680
rect 40498 256808 40554 256864
rect 40590 211928 40646 211984
rect 40498 45464 40554 45520
rect 40866 417968 40922 418024
rect 40774 408992 40830 409048
rect 41510 660320 41566 660376
rect 41694 660048 41750 660104
rect 41602 476720 41658 476776
rect 41050 387232 41106 387288
rect 40958 355952 41014 356008
rect 40958 50088 41014 50144
rect 59634 699896 59690 699952
rect 66258 699760 66314 699816
rect 73066 699896 73122 699952
rect 57794 666440 57850 666496
rect 55586 663992 55642 664048
rect 58806 663992 58862 664048
rect 73802 664264 73858 664320
rect 92938 700440 92994 700496
rect 116306 700576 116362 700632
rect 59910 662652 59966 662688
rect 59910 662632 59912 662652
rect 59912 662632 59964 662652
rect 59964 662632 59966 662652
rect 162858 700168 162914 700224
rect 59266 661952 59322 662008
rect 92386 661952 92442 662008
rect 229466 700984 229522 701040
rect 226154 700032 226210 700088
rect 240506 664400 240562 664456
rect 237470 664128 237526 664184
rect 255686 664264 255742 664320
rect 273902 664536 273958 664592
rect 295062 664672 295118 664728
rect 307206 663856 307262 663912
rect 322570 699896 322626 699952
rect 332690 699760 332746 699816
rect 349250 699760 349306 699816
rect 343638 668480 343694 668536
rect 346122 666440 346178 666496
rect 343454 664400 343510 664456
rect 349158 663720 349214 663776
rect 365994 699760 366050 699816
rect 399114 700848 399170 700904
rect 353298 662360 353354 662416
rect 284942 662088 284998 662144
rect 297822 662088 297878 662144
rect 301410 662088 301466 662144
rect 354034 662088 354090 662144
rect 358266 662088 358322 662144
rect 214654 661952 214710 662008
rect 243910 661952 243966 662008
rect 353022 661952 353078 662008
rect 166262 661816 166318 661872
rect 179510 661816 179566 661872
rect 192390 661816 192446 661872
rect 355966 661816 356022 661872
rect 367282 661816 367338 661872
rect 394790 661816 394846 661872
rect 449162 700712 449218 700768
rect 452474 700168 452530 700224
rect 437478 664264 437534 664320
rect 449346 663856 449402 663912
rect 469034 699760 469090 699816
rect 489090 699760 489146 699816
rect 502338 700848 502394 700904
rect 503994 664808 504050 664864
rect 440238 661816 440294 661872
rect 452106 661816 452162 661872
rect 461122 661816 461178 661872
rect 467194 661816 467250 661872
rect 512642 661680 512698 661736
rect 515218 661700 515274 661736
rect 528190 663856 528246 663912
rect 538954 699760 539010 699816
rect 528558 661816 528614 661872
rect 515218 661680 515220 661700
rect 515220 661680 515272 661700
rect 515272 661680 515274 661700
rect 524786 661680 524842 661736
rect 541898 661544 541954 661600
rect 542082 700304 542138 700360
rect 542082 660864 542138 660920
rect 541990 610816 542046 610872
rect 541990 471824 542046 471880
rect 541990 466248 542046 466304
rect 541990 442448 542046 442504
rect 542082 439048 542138 439104
rect 541990 438912 542046 438968
rect 542082 438096 542138 438152
rect 541898 193296 541954 193352
rect 41878 44240 41934 44296
rect 541990 143928 542046 143984
rect 59266 42336 59322 42392
rect 68006 42200 68062 42256
rect 60094 39752 60150 39808
rect 56506 3440 56562 3496
rect 157430 42064 157486 42120
rect 73250 3576 73306 3632
rect 84290 39480 84346 39536
rect 83186 6160 83242 6216
rect 96434 4800 96490 4856
rect 99746 5344 99802 5400
rect 116490 3712 116546 3768
rect 106370 3440 106426 3496
rect 132682 39888 132738 39944
rect 165986 39616 166042 39672
rect 175278 39616 175334 39672
rect 187606 10240 187662 10296
rect 223946 42336 224002 42392
rect 284022 42336 284078 42392
rect 371698 42336 371754 42392
rect 230110 42064 230166 42120
rect 213826 8880 213882 8936
rect 209594 5072 209650 5128
rect 202970 3984 203026 4040
rect 256974 39344 257030 39400
rect 246210 6296 246266 6352
rect 239586 5208 239642 5264
rect 249522 3984 249578 4040
rect 285678 40568 285734 40624
rect 287334 39480 287390 39536
rect 287702 33496 287758 33552
rect 308494 39888 308550 39944
rect 309506 6432 309562 6488
rect 302882 5480 302938 5536
rect 317510 39208 317566 39264
rect 348238 41384 348294 41440
rect 339498 3848 339554 3904
rect 353850 40296 353906 40352
rect 354954 40296 355010 40352
rect 350538 39072 350594 39128
rect 354586 35808 354642 35864
rect 354586 26288 354642 26344
rect 354586 26152 354642 26208
rect 354586 16632 354642 16688
rect 354586 16496 354642 16552
rect 354586 6976 354642 7032
rect 359370 3848 359426 3904
rect 378138 38664 378194 38720
rect 362682 3032 362738 3088
rect 405554 42336 405610 42392
rect 381082 40160 381138 40216
rect 390282 40024 390338 40080
rect 393318 40024 393374 40080
rect 392674 2896 392730 2952
rect 423678 39072 423734 39128
rect 432602 38800 432658 38856
rect 402794 2896 402850 2952
rect 419354 4936 419410 4992
rect 412730 3032 412786 3088
rect 425978 3032 426034 3088
rect 432602 3032 432658 3088
rect 439410 3168 439466 3224
rect 462962 39344 463018 39400
rect 471978 38936 472034 38992
rect 476026 4936 476082 4992
rect 459282 3032 459338 3088
rect 479338 3304 479394 3360
rect 488538 33768 488594 33824
rect 515954 3576 516010 3632
rect 519266 3848 519322 3904
rect 528558 33768 528614 33824
rect 542174 117272 542230 117328
rect 542082 95104 542138 95160
rect 542542 660456 542598 660512
rect 542726 641824 542782 641880
rect 542634 633392 542690 633448
rect 542634 615168 542690 615224
rect 542542 530032 542598 530088
rect 542542 524456 542598 524512
rect 542634 503376 542690 503432
rect 542726 484472 542782 484528
rect 542634 480256 542690 480312
rect 542910 350240 542966 350296
rect 543646 651072 543702 651128
rect 543646 596980 543648 597000
rect 543648 596980 543700 597000
rect 543700 596980 543702 597000
rect 543646 596944 543702 596980
rect 543278 422320 543334 422376
rect 543094 355136 543150 355192
rect 542910 305224 542966 305280
rect 542818 301824 542874 301880
rect 542818 291624 542874 291680
rect 543002 202136 543058 202192
rect 543094 198328 543150 198384
rect 543278 153448 543334 153504
rect 543186 140120 543242 140176
rect 544014 655152 544070 655208
rect 543922 458224 543978 458280
rect 543922 435684 543924 435704
rect 543924 435684 543976 435704
rect 543976 435684 543978 435704
rect 543922 435648 543978 435684
rect 543922 431332 543924 431352
rect 543924 431332 543976 431352
rect 543976 431332 543978 431352
rect 543922 431296 543978 431332
rect 544106 628088 544162 628144
rect 544014 426672 544070 426728
rect 543922 413208 543978 413264
rect 543830 252048 543886 252104
rect 543830 180548 543832 180568
rect 543832 180548 543884 180568
rect 543884 180548 543886 180568
rect 543830 180512 543886 180548
rect 543830 167220 543832 167240
rect 543832 167220 543884 167240
rect 543884 167220 543886 167240
rect 543830 167184 543886 167220
rect 543830 162424 543886 162480
rect 543830 150456 543886 150512
rect 543830 139440 543886 139496
rect 543830 131280 543886 131336
rect 543738 108976 543794 109032
rect 543738 104216 543794 104272
rect 543462 86264 543518 86320
rect 543830 81912 543886 81968
rect 543738 77288 543794 77344
rect 543830 68448 543886 68504
rect 543830 64132 543832 64152
rect 543832 64132 543884 64152
rect 543884 64132 543886 64152
rect 543830 64096 543886 64132
rect 543830 59508 543832 59528
rect 543832 59508 543884 59528
rect 543884 59508 543886 59528
rect 543830 59472 543886 59508
rect 543830 54984 543886 55040
rect 543830 50632 543886 50688
rect 544014 372952 544070 373008
rect 544290 661408 544346 661464
rect 544198 475904 544254 475960
rect 544198 417732 544200 417752
rect 544200 417732 544252 417752
rect 544252 417732 544254 417752
rect 544198 417696 544254 417732
rect 544198 408720 544254 408776
rect 544198 381928 544254 381984
rect 544106 369144 544162 369200
rect 544106 368464 544162 368520
rect 544658 659504 544714 659560
rect 544658 547576 544714 547632
rect 544658 534112 544714 534168
rect 544658 520820 544660 520840
rect 544660 520820 544712 520840
rect 544712 520820 544714 520840
rect 544658 520784 544714 520820
rect 544658 511844 544660 511864
rect 544660 511844 544712 511864
rect 544712 511844 544714 511864
rect 544658 511808 544714 511844
rect 544658 507320 544714 507376
rect 544658 493892 544660 493912
rect 544660 493892 544712 493912
rect 544712 493892 544714 493912
rect 544658 493856 544714 493892
rect 544658 489540 544660 489560
rect 544660 489540 544712 489560
rect 544712 489540 544714 489560
rect 544658 489504 544714 489540
rect 544658 466792 544714 466848
rect 544658 462612 544660 462632
rect 544660 462612 544712 462632
rect 544712 462612 544714 462632
rect 544658 462576 544714 462612
rect 544658 453464 544714 453520
rect 544658 449248 544714 449304
rect 544658 445712 544714 445768
rect 544566 346160 544622 346216
rect 544566 337048 544622 337104
rect 544474 332832 544530 332888
rect 544382 328208 544438 328264
rect 544290 323856 544346 323912
rect 544290 314744 544346 314800
rect 544382 310120 544438 310176
rect 544474 229780 544476 229800
rect 544476 229780 544528 229800
rect 544528 229780 544530 229800
rect 544474 229744 544530 229780
rect 544474 211656 544530 211712
rect 544474 191664 544530 191720
rect 544474 171400 544530 171456
rect 544474 122168 544530 122224
rect 544842 646176 544898 646232
rect 544842 637200 544898 637256
rect 544842 623872 544898 623928
rect 544842 619112 544898 619168
rect 544842 605956 544844 605976
rect 544844 605956 544896 605976
rect 544896 605956 544898 605976
rect 544842 605920 544898 605956
rect 544842 601160 544898 601216
rect 544934 574676 544936 574696
rect 544936 574676 544988 574696
rect 544988 574676 544990 574696
rect 544934 574640 544990 574676
rect 544934 570016 544990 570072
rect 544934 565664 544990 565720
rect 545026 561040 545082 561096
rect 544934 552100 544936 552120
rect 544936 552100 544988 552120
rect 544988 552100 544990 552120
rect 544934 552064 544990 552100
rect 544934 538736 544990 538792
rect 545026 516296 545082 516352
rect 545026 498344 545082 498400
rect 544934 440308 544936 440328
rect 544936 440308 544988 440328
rect 544988 440308 544990 440328
rect 544934 440272 544990 440308
rect 544934 404368 544990 404424
rect 544750 400016 544806 400072
rect 544750 395392 544806 395448
rect 544750 390904 544806 390960
rect 544750 377476 544752 377496
rect 544752 377476 544804 377496
rect 544804 377476 544806 377496
rect 544750 377440 544806 377476
rect 544750 364148 544752 364168
rect 544752 364148 544804 364168
rect 544804 364148 544806 364168
rect 544750 364112 544806 364148
rect 544934 386416 544990 386472
rect 544934 359352 544990 359408
rect 544750 341808 544806 341864
rect 544934 319096 544990 319152
rect 544934 278840 544990 278896
rect 544750 274624 544806 274680
rect 544934 269864 544990 269920
rect 544750 256536 544806 256592
rect 544750 247560 544806 247616
rect 544750 242956 544806 242992
rect 544750 242936 544752 242956
rect 544752 242936 544804 242956
rect 544804 242936 544806 242956
rect 544750 238584 544806 238640
rect 544750 225256 544806 225312
rect 544750 220632 544806 220688
rect 544750 207440 544806 207496
rect 544750 184728 544806 184784
rect 544750 175888 544806 175944
rect 544750 158208 544806 158264
rect 544658 149232 544714 149288
rect 544658 113328 544714 113384
rect 544658 99864 544714 99920
rect 544750 90888 544806 90944
rect 544658 46144 544714 46200
rect 545026 126520 545082 126576
rect 545302 578312 545358 578368
rect 545302 556552 545358 556608
rect 545670 287816 545726 287872
rect 545486 265512 545542 265568
rect 545578 216280 545634 216336
rect 545670 189352 545726 189408
rect 545670 72936 545726 72992
rect 547050 291080 547106 291136
rect 550822 482160 550878 482216
rect 551650 39616 551706 39672
rect 552662 663992 552718 664048
rect 552018 44104 552074 44160
rect 562322 653384 562378 653440
rect 554778 43560 554834 43616
rect 580630 696360 580686 696416
rect 580170 691464 580226 691520
rect 579618 686568 579674 686624
rect 580170 681672 580226 681728
rect 580170 671880 580226 671936
rect 579618 666984 579674 667040
rect 579618 662088 579674 662144
rect 580078 642232 580134 642288
rect 579986 637336 580042 637392
rect 580170 632440 580226 632496
rect 580170 622648 580226 622704
rect 579986 617752 580042 617808
rect 579618 612856 579674 612912
rect 580170 607960 580226 608016
rect 579618 603064 579674 603120
rect 580170 598168 580226 598224
rect 579618 593000 579674 593056
rect 580170 588104 580226 588160
rect 579986 583208 580042 583264
rect 579618 578312 579674 578368
rect 580170 573416 580226 573472
rect 580170 558728 580226 558784
rect 580170 553832 580226 553888
rect 580078 544040 580134 544096
rect 580170 538872 580226 538928
rect 580262 533976 580318 534032
rect 580170 529080 580226 529136
rect 579618 524184 579674 524240
rect 580262 519288 580318 519344
rect 580170 514392 580226 514448
rect 579986 504600 580042 504656
rect 579710 499704 579766 499760
rect 579986 494808 580042 494864
rect 580170 489932 580226 489968
rect 580170 489912 580172 489932
rect 580172 489912 580224 489932
rect 580224 489912 580226 489932
rect 580170 484744 580226 484800
rect 579618 479848 579674 479904
rect 580170 474952 580226 475008
rect 579986 470056 580042 470112
rect 580170 460264 580226 460320
rect 580170 455368 580226 455424
rect 580170 450472 580226 450528
rect 580170 445576 580226 445632
rect 580170 440680 580226 440736
rect 580170 435784 580226 435840
rect 579618 430616 579674 430672
rect 580170 425720 580226 425776
rect 580170 411032 580226 411088
rect 580170 406136 580226 406192
rect 579710 401240 579766 401296
rect 579618 391448 579674 391504
rect 580170 386552 580226 386608
rect 579802 381656 579858 381712
rect 580170 376488 580226 376544
rect 579618 371592 579674 371648
rect 580170 366696 580226 366752
rect 580170 361800 580226 361856
rect 579986 356904 580042 356960
rect 580170 352008 580226 352064
rect 580170 347112 580226 347168
rect 580170 337320 580226 337376
rect 579986 327528 580042 327584
rect 579802 322360 579858 322416
rect 580170 312568 580226 312624
rect 580170 307708 580172 307728
rect 580172 307708 580224 307728
rect 580224 307708 580226 307728
rect 580170 307672 580226 307708
rect 580170 302776 580226 302832
rect 579618 297880 579674 297936
rect 579802 292984 579858 293040
rect 579618 288088 579674 288144
rect 579618 283192 579674 283248
rect 579986 278296 580042 278352
rect 580170 273400 580226 273456
rect 580170 258440 580226 258496
rect 579802 253544 579858 253600
rect 579618 248648 579674 248704
rect 580170 238856 580226 238912
rect 579986 233960 580042 234016
rect 580170 229100 580172 229120
rect 580172 229100 580224 229120
rect 580224 229100 580226 229120
rect 580170 229064 580226 229100
rect 579802 219272 579858 219328
rect 580170 214104 580226 214160
rect 579986 209208 580042 209264
rect 580170 199416 580226 199472
rect 580170 194540 580226 194576
rect 580170 194520 580172 194540
rect 580172 194520 580224 194540
rect 580224 194520 580226 194540
rect 579618 189624 579674 189680
rect 580170 184728 580226 184784
rect 579986 179832 580042 179888
rect 579618 174936 579674 174992
rect 579986 165144 580042 165200
rect 580170 160012 580172 160032
rect 580172 160012 580224 160032
rect 580224 160012 580226 160032
rect 580170 159976 580226 160012
rect 579618 155080 579674 155136
rect 579618 150184 579674 150240
rect 580170 140392 580226 140448
rect 579618 135496 579674 135552
rect 579802 130600 579858 130656
rect 580170 120808 580226 120864
rect 579618 115912 579674 115968
rect 580170 111016 580226 111072
rect 580170 105848 580226 105904
rect 579618 100952 579674 101008
rect 578974 96056 579030 96112
rect 578882 86264 578938 86320
rect 580170 81388 580226 81424
rect 580170 81368 580172 81388
rect 580172 81368 580224 81388
rect 580224 81368 580226 81388
rect 580170 61784 580226 61840
rect 580078 56888 580134 56944
rect 579986 51720 580042 51776
rect 579986 46860 579988 46880
rect 579988 46860 580040 46880
rect 580040 46860 580042 46880
rect 579986 46824 580042 46860
rect 580170 41928 580226 41984
rect 580906 676776 580962 676832
rect 580630 652296 580686 652352
rect 580538 548936 580594 548992
rect 580538 509496 580594 509552
rect 580538 465160 580594 465216
rect 580630 420824 580686 420880
rect 580538 415928 580594 415984
rect 580446 268232 580502 268288
rect 580446 263336 580502 263392
rect 580354 243752 580410 243808
rect 580354 204312 580410 204368
rect 580630 396344 580686 396400
rect 580814 657192 580870 657248
rect 580722 342216 580778 342272
rect 580722 332424 580778 332480
rect 580814 317464 580870 317520
rect 580906 170040 580962 170096
rect 580722 125704 580778 125760
rect 580814 71576 580870 71632
rect 580170 37032 580226 37088
rect 580078 32136 580134 32192
rect 580078 27240 580134 27296
rect 580722 44648 580778 44704
rect 580446 22344 580502 22400
rect 580906 66680 580962 66736
rect 580722 12552 580778 12608
rect 580170 7656 580226 7712
rect 580170 2760 580226 2816
<< metal3 >>
rect -960 703762 480 703852
rect 3417 703762 3483 703765
rect -960 703760 3483 703762
rect -960 703704 3422 703760
rect 3478 703704 3483 703760
rect -960 703702 3483 703704
rect -960 703612 480 703702
rect 3417 703699 3483 703702
rect 583520 701164 584960 701404
rect 229461 701042 229527 701045
rect 541934 701042 541940 701044
rect 229461 701040 541940 701042
rect 229461 700984 229466 701040
rect 229522 700984 541940 701040
rect 229461 700982 541940 700984
rect 229461 700979 229527 700982
rect 541934 700980 541940 700982
rect 542004 700980 542010 701044
rect 39614 700844 39620 700908
rect 39684 700906 39690 700908
rect 399109 700906 399175 700909
rect 39684 700904 399175 700906
rect 39684 700848 399114 700904
rect 399170 700848 399175 700904
rect 39684 700846 399175 700848
rect 39684 700844 39690 700846
rect 399109 700843 399175 700846
rect 405590 700844 405596 700908
rect 405660 700906 405666 700908
rect 502333 700906 502399 700909
rect 405660 700904 502399 700906
rect 405660 700848 502338 700904
rect 502394 700848 502399 700904
rect 405660 700846 502399 700848
rect 405660 700844 405666 700846
rect 502333 700843 502399 700846
rect 39062 700708 39068 700772
rect 39132 700770 39138 700772
rect 449157 700770 449223 700773
rect 39132 700768 449223 700770
rect 39132 700712 449162 700768
rect 449218 700712 449223 700768
rect 39132 700710 449223 700712
rect 39132 700708 39138 700710
rect 449157 700707 449223 700710
rect 116301 700634 116367 700637
rect 542854 700634 542860 700636
rect 116301 700632 542860 700634
rect 116301 700576 116306 700632
rect 116362 700576 542860 700632
rect 116301 700574 542860 700576
rect 116301 700571 116367 700574
rect 542854 700572 542860 700574
rect 542924 700572 542930 700636
rect 92933 700498 92999 700501
rect 542486 700498 542492 700500
rect 92933 700496 542492 700498
rect 92933 700440 92938 700496
rect 92994 700440 542492 700496
rect 92933 700438 542492 700440
rect 92933 700435 92999 700438
rect 542486 700436 542492 700438
rect 542556 700436 542562 700500
rect 40534 700300 40540 700364
rect 40604 700362 40610 700364
rect 542077 700362 542143 700365
rect 40604 700360 542143 700362
rect 40604 700304 542082 700360
rect 542138 700304 542143 700360
rect 40604 700302 542143 700304
rect 40604 700300 40610 700302
rect 542077 700299 542143 700302
rect 162853 700226 162919 700229
rect 370446 700226 370452 700228
rect 162853 700224 370452 700226
rect 162853 700168 162858 700224
rect 162914 700168 370452 700224
rect 162853 700166 370452 700168
rect 162853 700163 162919 700166
rect 370446 700164 370452 700166
rect 370516 700164 370522 700228
rect 415894 700164 415900 700228
rect 415964 700226 415970 700228
rect 452469 700226 452535 700229
rect 415964 700224 452535 700226
rect 415964 700168 452474 700224
rect 452530 700168 452535 700224
rect 415964 700166 452535 700168
rect 415964 700164 415970 700166
rect 452469 700163 452535 700166
rect 226149 700090 226215 700093
rect 362166 700090 362172 700092
rect 226149 700088 362172 700090
rect 226149 700032 226154 700088
rect 226210 700032 362172 700088
rect 226149 700030 362172 700032
rect 226149 700027 226215 700030
rect 362166 700028 362172 700030
rect 362236 700028 362242 700092
rect 59629 699954 59695 699957
rect 59854 699954 59860 699956
rect 59629 699952 59860 699954
rect 59629 699896 59634 699952
rect 59690 699896 59860 699952
rect 59629 699894 59860 699896
rect 59629 699891 59695 699894
rect 59854 699892 59860 699894
rect 59924 699892 59930 699956
rect 73061 699954 73127 699957
rect 64830 699952 73127 699954
rect 64830 699896 73066 699952
rect 73122 699896 73127 699952
rect 64830 699894 73127 699896
rect 39982 699756 39988 699820
rect 40052 699818 40058 699820
rect 64830 699818 64890 699894
rect 73061 699891 73127 699894
rect 322565 699954 322631 699957
rect 364926 699954 364932 699956
rect 322565 699952 364932 699954
rect 322565 699896 322570 699952
rect 322626 699896 364932 699952
rect 322565 699894 364932 699896
rect 322565 699891 322631 699894
rect 364926 699892 364932 699894
rect 364996 699892 365002 699956
rect 367686 699954 367692 699956
rect 365486 699894 367692 699954
rect 66253 699820 66319 699821
rect 66253 699818 66300 699820
rect 40052 699758 64890 699818
rect 66208 699816 66300 699818
rect 66208 699760 66258 699816
rect 66208 699758 66300 699760
rect 40052 699756 40058 699758
rect 66253 699756 66300 699758
rect 66364 699756 66370 699820
rect 332685 699818 332751 699821
rect 333830 699818 333836 699820
rect 332685 699816 333836 699818
rect 332685 699760 332690 699816
rect 332746 699760 333836 699816
rect 332685 699758 333836 699760
rect 66253 699755 66319 699756
rect 332685 699755 332751 699758
rect 333830 699756 333836 699758
rect 333900 699756 333906 699820
rect 349245 699818 349311 699821
rect 365486 699818 365546 699894
rect 367686 699892 367692 699894
rect 367756 699892 367762 699956
rect 349245 699816 365546 699818
rect 349245 699760 349250 699816
rect 349306 699760 365546 699816
rect 349245 699758 365546 699760
rect 349245 699755 349311 699758
rect 365662 699756 365668 699820
rect 365732 699818 365738 699820
rect 365989 699818 366055 699821
rect 365732 699816 366055 699818
rect 365732 699760 365994 699816
rect 366050 699760 366055 699816
rect 365732 699758 366055 699760
rect 365732 699756 365738 699758
rect 365989 699755 366055 699758
rect 467782 699756 467788 699820
rect 467852 699818 467858 699820
rect 469029 699818 469095 699821
rect 467852 699816 469095 699818
rect 467852 699760 469034 699816
rect 469090 699760 469095 699816
rect 467852 699758 469095 699760
rect 467852 699756 467858 699758
rect 469029 699755 469095 699758
rect 488574 699756 488580 699820
rect 488644 699818 488650 699820
rect 489085 699818 489151 699821
rect 488644 699816 489151 699818
rect 488644 699760 489090 699816
rect 489146 699760 489151 699816
rect 488644 699758 489151 699760
rect 488644 699756 488650 699758
rect 489085 699755 489151 699758
rect 538949 699818 539015 699821
rect 543774 699818 543780 699820
rect 538949 699816 543780 699818
rect 538949 699760 538954 699816
rect 539010 699760 543780 699816
rect 538949 699758 543780 699760
rect 538949 699755 539015 699758
rect 543774 699756 543780 699758
rect 543844 699756 543850 699820
rect -960 698594 480 698684
rect 3233 698594 3299 698597
rect -960 698592 3299 698594
rect -960 698536 3238 698592
rect 3294 698536 3299 698592
rect -960 698534 3299 698536
rect -960 698444 480 698534
rect 3233 698531 3299 698534
rect 580625 696418 580691 696421
rect 583520 696418 584960 696508
rect 580625 696416 584960 696418
rect 580625 696360 580630 696416
rect 580686 696360 584960 696416
rect 580625 696358 584960 696360
rect 580625 696355 580691 696358
rect 583520 696268 584960 696358
rect -960 693698 480 693788
rect 3141 693698 3207 693701
rect -960 693696 3207 693698
rect -960 693640 3146 693696
rect 3202 693640 3207 693696
rect -960 693638 3207 693640
rect -960 693548 480 693638
rect 3141 693635 3207 693638
rect 580165 691522 580231 691525
rect 583520 691522 584960 691612
rect 580165 691520 584960 691522
rect 580165 691464 580170 691520
rect 580226 691464 584960 691520
rect 580165 691462 584960 691464
rect 580165 691459 580231 691462
rect 583520 691372 584960 691462
rect -960 688802 480 688892
rect 3509 688802 3575 688805
rect -960 688800 3575 688802
rect -960 688744 3514 688800
rect 3570 688744 3575 688800
rect -960 688742 3575 688744
rect -960 688652 480 688742
rect 3509 688739 3575 688742
rect 579613 686626 579679 686629
rect 583520 686626 584960 686716
rect 579613 686624 584960 686626
rect 579613 686568 579618 686624
rect 579674 686568 584960 686624
rect 579613 686566 584960 686568
rect 579613 686563 579679 686566
rect 583520 686476 584960 686566
rect -960 683906 480 683996
rect 3417 683906 3483 683909
rect -960 683904 3483 683906
rect -960 683848 3422 683904
rect 3478 683848 3483 683904
rect -960 683846 3483 683848
rect -960 683756 480 683846
rect 3417 683843 3483 683846
rect 580165 681730 580231 681733
rect 583520 681730 584960 681820
rect 580165 681728 584960 681730
rect 580165 681672 580170 681728
rect 580226 681672 584960 681728
rect 580165 681670 584960 681672
rect 580165 681667 580231 681670
rect 583520 681580 584960 681670
rect -960 679010 480 679100
rect 3877 679010 3943 679013
rect -960 679008 3943 679010
rect -960 678952 3882 679008
rect 3938 678952 3943 679008
rect -960 678950 3943 678952
rect -960 678860 480 678950
rect 3877 678947 3943 678950
rect 580901 676834 580967 676837
rect 583520 676834 584960 676924
rect 580901 676832 584960 676834
rect 580901 676776 580906 676832
rect 580962 676776 584960 676832
rect 580901 676774 584960 676776
rect 580901 676771 580967 676774
rect 583520 676684 584960 676774
rect -960 674114 480 674204
rect 3693 674114 3759 674117
rect -960 674112 3759 674114
rect -960 674056 3698 674112
rect 3754 674056 3759 674112
rect -960 674054 3759 674056
rect -960 673964 480 674054
rect 3693 674051 3759 674054
rect 580165 671938 580231 671941
rect 583520 671938 584960 672028
rect 580165 671936 584960 671938
rect 580165 671880 580170 671936
rect 580226 671880 584960 671936
rect 580165 671878 584960 671880
rect 580165 671875 580231 671878
rect 583520 671788 584960 671878
rect -960 669218 480 669308
rect 3785 669218 3851 669221
rect -960 669216 3851 669218
rect -960 669160 3790 669216
rect 3846 669160 3851 669216
rect -960 669158 3851 669160
rect -960 669068 480 669158
rect 3785 669155 3851 669158
rect 343633 668538 343699 668541
rect 353334 668538 353340 668540
rect 343633 668536 353340 668538
rect 343633 668480 343638 668536
rect 343694 668480 353340 668536
rect 343633 668478 353340 668480
rect 343633 668475 343699 668478
rect 353334 668476 353340 668478
rect 353404 668476 353410 668540
rect 579613 667042 579679 667045
rect 583520 667042 584960 667132
rect 579613 667040 584960 667042
rect 579613 666984 579618 667040
rect 579674 666984 584960 667040
rect 579613 666982 584960 666984
rect 579613 666979 579679 666982
rect 583520 666892 584960 666982
rect 55990 666436 55996 666500
rect 56060 666498 56066 666500
rect 57789 666498 57855 666501
rect 56060 666496 57855 666498
rect 56060 666440 57794 666496
rect 57850 666440 57855 666496
rect 56060 666438 57855 666440
rect 56060 666436 56066 666438
rect 57789 666435 57855 666438
rect 346117 666498 346183 666501
rect 351862 666498 351868 666500
rect 346117 666496 351868 666498
rect 346117 666440 346122 666496
rect 346178 666440 351868 666496
rect 346117 666438 351868 666440
rect 346117 666435 346183 666438
rect 351862 666436 351868 666438
rect 351932 666436 351938 666500
rect 8937 664866 9003 664869
rect 503989 664866 504055 664869
rect 8937 664864 504055 664866
rect 8937 664808 8942 664864
rect 8998 664808 503994 664864
rect 504050 664808 504055 664864
rect 8937 664806 504055 664808
rect 8937 664803 9003 664806
rect 503989 664803 504055 664806
rect 295057 664730 295123 664733
rect 368974 664730 368980 664732
rect 295057 664728 368980 664730
rect 295057 664672 295062 664728
rect 295118 664672 368980 664728
rect 295057 664670 368980 664672
rect 295057 664667 295123 664670
rect 368974 664668 368980 664670
rect 369044 664668 369050 664732
rect 273897 664594 273963 664597
rect 363454 664594 363460 664596
rect 273897 664592 363460 664594
rect 273897 664536 273902 664592
rect 273958 664536 363460 664592
rect 273897 664534 363460 664536
rect 273897 664531 273963 664534
rect 363454 664532 363460 664534
rect 363524 664532 363530 664596
rect -960 664322 480 664412
rect 42742 664396 42748 664460
rect 42812 664458 42818 664460
rect 240501 664458 240567 664461
rect 42812 664456 240567 664458
rect 42812 664400 240506 664456
rect 240562 664400 240567 664456
rect 42812 664398 240567 664400
rect 42812 664396 42818 664398
rect 240501 664395 240567 664398
rect 343449 664458 343515 664461
rect 436686 664458 436692 664460
rect 343449 664456 436692 664458
rect 343449 664400 343454 664456
rect 343510 664400 436692 664456
rect 343449 664398 436692 664400
rect 343449 664395 343515 664398
rect 436686 664396 436692 664398
rect 436756 664396 436762 664460
rect 3417 664322 3483 664325
rect -960 664320 3483 664322
rect -960 664264 3422 664320
rect 3478 664264 3483 664320
rect -960 664262 3483 664264
rect -960 664172 480 664262
rect 3417 664259 3483 664262
rect 55070 664260 55076 664324
rect 55140 664322 55146 664324
rect 73797 664322 73863 664325
rect 55140 664320 73863 664322
rect 55140 664264 73802 664320
rect 73858 664264 73863 664320
rect 55140 664262 73863 664264
rect 55140 664260 55146 664262
rect 73797 664259 73863 664262
rect 255681 664322 255747 664325
rect 360694 664322 360700 664324
rect 255681 664320 360700 664322
rect 255681 664264 255686 664320
rect 255742 664264 360700 664320
rect 255681 664262 360700 664264
rect 255681 664259 255747 664262
rect 360694 664260 360700 664262
rect 360764 664260 360770 664324
rect 402830 664260 402836 664324
rect 402900 664322 402906 664324
rect 437473 664322 437539 664325
rect 402900 664320 437539 664322
rect 402900 664264 437478 664320
rect 437534 664264 437539 664320
rect 402900 664262 437539 664264
rect 402900 664260 402906 664262
rect 437473 664259 437539 664262
rect 237465 664186 237531 664189
rect 545062 664186 545068 664188
rect 237465 664184 545068 664186
rect 237465 664128 237470 664184
rect 237526 664128 545068 664184
rect 237465 664126 545068 664128
rect 237465 664123 237531 664126
rect 545062 664124 545068 664126
rect 545132 664124 545138 664188
rect 42374 663988 42380 664052
rect 42444 664050 42450 664052
rect 55581 664050 55647 664053
rect 42444 664048 55647 664050
rect 42444 663992 55586 664048
rect 55642 663992 55647 664048
rect 42444 663990 55647 663992
rect 42444 663988 42450 663990
rect 55581 663987 55647 663990
rect 58801 664050 58867 664053
rect 552657 664050 552723 664053
rect 58801 664048 552723 664050
rect 58801 663992 58806 664048
rect 58862 663992 552662 664048
rect 552718 663992 552723 664048
rect 58801 663990 552723 663992
rect 58801 663987 58867 663990
rect 552657 663987 552723 663990
rect 307201 663914 307267 663917
rect 310462 663914 310468 663916
rect 307201 663912 310468 663914
rect 307201 663856 307206 663912
rect 307262 663856 310468 663912
rect 307201 663854 310468 663856
rect 307201 663851 307267 663854
rect 310462 663852 310468 663854
rect 310532 663852 310538 663916
rect 443494 663852 443500 663916
rect 443564 663914 443570 663916
rect 449341 663914 449407 663917
rect 443564 663912 449407 663914
rect 443564 663856 449346 663912
rect 449402 663856 449407 663912
rect 443564 663854 449407 663856
rect 443564 663852 443570 663854
rect 449341 663851 449407 663854
rect 528185 663914 528251 663917
rect 541014 663914 541020 663916
rect 528185 663912 541020 663914
rect 528185 663856 528190 663912
rect 528246 663856 541020 663912
rect 528185 663854 541020 663856
rect 528185 663851 528251 663854
rect 541014 663852 541020 663854
rect 541084 663852 541090 663916
rect 349153 663778 349219 663781
rect 354806 663778 354812 663780
rect 349153 663776 354812 663778
rect 349153 663720 349158 663776
rect 349214 663720 354812 663776
rect 349153 663718 354812 663720
rect 349153 663715 349219 663718
rect 354806 663716 354812 663718
rect 354876 663716 354882 663780
rect 59905 662692 59971 662693
rect 59854 662690 59860 662692
rect 59814 662630 59860 662690
rect 59924 662688 59971 662692
rect 59966 662632 59971 662688
rect 59854 662628 59860 662630
rect 59924 662628 59971 662632
rect 59905 662627 59971 662628
rect 353293 662418 353359 662421
rect 355358 662418 355364 662420
rect 353293 662416 355364 662418
rect 353293 662360 353298 662416
rect 353354 662360 355364 662416
rect 353293 662358 355364 662360
rect 353293 662355 353359 662358
rect 355358 662356 355364 662358
rect 355428 662356 355434 662420
rect 356094 662282 356100 662284
rect 335310 662222 356100 662282
rect 284937 662146 285003 662149
rect 285806 662146 285812 662148
rect 284937 662144 285812 662146
rect 284937 662088 284942 662144
rect 284998 662088 285812 662144
rect 284937 662086 285812 662088
rect 284937 662083 285003 662086
rect 285806 662084 285812 662086
rect 285876 662084 285882 662148
rect 297817 662146 297883 662149
rect 301405 662148 301471 662149
rect 297950 662146 297956 662148
rect 297817 662144 297956 662146
rect 297817 662088 297822 662144
rect 297878 662088 297956 662144
rect 297817 662086 297956 662088
rect 297817 662083 297883 662086
rect 297950 662084 297956 662086
rect 298020 662084 298026 662148
rect 301405 662144 301452 662148
rect 301516 662146 301522 662148
rect 301405 662088 301410 662144
rect 301405 662084 301452 662088
rect 301516 662086 301562 662146
rect 301516 662084 301522 662086
rect 301405 662083 301471 662084
rect 53230 661948 53236 662012
rect 53300 662010 53306 662012
rect 59261 662010 59327 662013
rect 53300 662008 59327 662010
rect 53300 661952 59266 662008
rect 59322 661952 59327 662008
rect 53300 661950 59327 661952
rect 53300 661948 53306 661950
rect 59261 661947 59327 661950
rect 92381 662010 92447 662013
rect 98678 662010 98684 662012
rect 92381 662008 98684 662010
rect 92381 661952 92386 662008
rect 92442 661952 98684 662008
rect 92381 661950 98684 661952
rect 92381 661947 92447 661950
rect 98678 661948 98684 661950
rect 98748 661948 98754 662012
rect 172462 661948 172468 662012
rect 172532 662010 172538 662012
rect 214649 662010 214715 662013
rect 172532 662008 214715 662010
rect 172532 661952 214654 662008
rect 214710 661952 214715 662008
rect 172532 661950 214715 661952
rect 172532 661948 172538 661950
rect 214649 661947 214715 661950
rect 243905 662010 243971 662013
rect 335310 662010 335370 662222
rect 356094 662220 356100 662222
rect 356164 662220 356170 662284
rect 354029 662148 354095 662149
rect 354029 662146 354076 662148
rect 353984 662144 354076 662146
rect 353984 662088 354034 662144
rect 353984 662086 354076 662088
rect 354029 662084 354076 662086
rect 354140 662084 354146 662148
rect 358261 662146 358327 662149
rect 358670 662146 358676 662148
rect 358261 662144 358676 662146
rect 358261 662088 358266 662144
rect 358322 662088 358676 662144
rect 358261 662086 358676 662088
rect 354029 662083 354095 662084
rect 358261 662083 358327 662086
rect 358670 662084 358676 662086
rect 358740 662084 358746 662148
rect 579613 662146 579679 662149
rect 583520 662146 584960 662236
rect 579613 662144 584960 662146
rect 579613 662088 579618 662144
rect 579674 662088 584960 662144
rect 579613 662086 584960 662088
rect 579613 662083 579679 662086
rect 243905 662008 335370 662010
rect 243905 661952 243910 662008
rect 243966 661952 335370 662008
rect 243905 661950 335370 661952
rect 353017 662010 353083 662013
rect 354438 662010 354444 662012
rect 353017 662008 354444 662010
rect 353017 661952 353022 662008
rect 353078 661952 354444 662008
rect 353017 661950 354444 661952
rect 243905 661947 243971 661950
rect 353017 661947 353083 661950
rect 354438 661948 354444 661950
rect 354508 661948 354514 662012
rect 358854 662010 358860 662012
rect 354630 661950 358860 662010
rect 53414 661812 53420 661876
rect 53484 661874 53490 661876
rect 166257 661874 166323 661877
rect 179505 661876 179571 661877
rect 179454 661874 179460 661876
rect 53484 661872 166323 661874
rect 53484 661816 166262 661872
rect 166318 661816 166323 661872
rect 53484 661814 166323 661816
rect 179414 661814 179460 661874
rect 179524 661872 179571 661876
rect 179566 661816 179571 661872
rect 53484 661812 53490 661814
rect 166257 661811 166323 661814
rect 179454 661812 179460 661814
rect 179524 661812 179571 661816
rect 179505 661811 179571 661812
rect 192385 661874 192451 661877
rect 354630 661874 354690 661950
rect 358854 661948 358860 661950
rect 358924 661948 358930 662012
rect 583520 661996 584960 662086
rect 192385 661872 354690 661874
rect 192385 661816 192390 661872
rect 192446 661816 354690 661872
rect 192385 661814 354690 661816
rect 355961 661874 356027 661877
rect 356646 661874 356652 661876
rect 355961 661872 356652 661874
rect 355961 661816 355966 661872
rect 356022 661816 356652 661872
rect 355961 661814 356652 661816
rect 192385 661811 192451 661814
rect 355961 661811 356027 661814
rect 356646 661812 356652 661814
rect 356716 661812 356722 661876
rect 366030 661812 366036 661876
rect 366100 661874 366106 661876
rect 367277 661874 367343 661877
rect 394785 661876 394851 661877
rect 440233 661876 440299 661877
rect 394734 661874 394740 661876
rect 366100 661872 367343 661874
rect 366100 661816 367282 661872
rect 367338 661816 367343 661872
rect 366100 661814 367343 661816
rect 394694 661814 394740 661874
rect 394804 661872 394851 661876
rect 440182 661874 440188 661876
rect 394846 661816 394851 661872
rect 366100 661812 366106 661814
rect 367277 661811 367343 661814
rect 394734 661812 394740 661814
rect 394804 661812 394851 661816
rect 440142 661814 440188 661874
rect 440252 661872 440299 661876
rect 440294 661816 440299 661872
rect 440182 661812 440188 661814
rect 440252 661812 440299 661816
rect 451038 661812 451044 661876
rect 451108 661874 451114 661876
rect 452101 661874 452167 661877
rect 451108 661872 452167 661874
rect 451108 661816 452106 661872
rect 452162 661816 452167 661872
rect 451108 661814 452167 661816
rect 451108 661812 451114 661814
rect 394785 661811 394851 661812
rect 440233 661811 440299 661812
rect 452101 661811 452167 661814
rect 460974 661812 460980 661876
rect 461044 661874 461050 661876
rect 461117 661874 461183 661877
rect 461044 661872 461183 661874
rect 461044 661816 461122 661872
rect 461178 661816 461183 661872
rect 461044 661814 461183 661816
rect 461044 661812 461050 661814
rect 461117 661811 461183 661814
rect 466494 661812 466500 661876
rect 466564 661874 466570 661876
rect 467189 661874 467255 661877
rect 528553 661874 528619 661877
rect 466564 661872 467255 661874
rect 466564 661816 467194 661872
rect 467250 661816 467255 661872
rect 466564 661814 467255 661816
rect 466564 661812 466570 661814
rect 467189 661811 467255 661814
rect 509190 661872 528619 661874
rect 509190 661816 528558 661872
rect 528614 661816 528619 661872
rect 509190 661814 528619 661816
rect 38878 661676 38884 661740
rect 38948 661738 38954 661740
rect 509190 661738 509250 661814
rect 528553 661811 528619 661814
rect 38948 661678 509250 661738
rect 38948 661676 38954 661678
rect 512126 661676 512132 661740
rect 512196 661738 512202 661740
rect 512637 661738 512703 661741
rect 515213 661740 515279 661741
rect 515213 661738 515260 661740
rect 512196 661736 512703 661738
rect 512196 661680 512642 661736
rect 512698 661680 512703 661736
rect 512196 661678 512703 661680
rect 515168 661736 515260 661738
rect 515168 661680 515218 661736
rect 515168 661678 515260 661680
rect 512196 661676 512202 661678
rect 512637 661675 512703 661678
rect 515213 661676 515260 661678
rect 515324 661676 515330 661740
rect 524454 661676 524460 661740
rect 524524 661738 524530 661740
rect 524781 661738 524847 661741
rect 524524 661736 524847 661738
rect 524524 661680 524786 661736
rect 524842 661680 524847 661736
rect 524524 661678 524847 661680
rect 524524 661676 524530 661678
rect 515213 661675 515279 661676
rect 524781 661675 524847 661678
rect 121494 661540 121500 661604
rect 121564 661602 121570 661604
rect 541893 661602 541959 661605
rect 121564 661600 541959 661602
rect 121564 661544 541898 661600
rect 541954 661544 541959 661600
rect 121564 661542 541959 661544
rect 121564 661540 121570 661542
rect 541893 661539 541959 661542
rect 108982 661404 108988 661468
rect 109052 661466 109058 661468
rect 544285 661466 544351 661469
rect 109052 661464 544351 661466
rect 109052 661408 544290 661464
rect 544346 661408 544351 661464
rect 109052 661406 544351 661408
rect 109052 661404 109058 661406
rect 544285 661403 544351 661406
rect 49734 661268 49740 661332
rect 49804 661330 49810 661332
rect 541750 661330 541756 661332
rect 49804 661270 541756 661330
rect 49804 661268 49810 661270
rect 541750 661268 541756 661270
rect 541820 661268 541826 661332
rect 6269 661194 6335 661197
rect 366030 661194 366036 661196
rect 6269 661192 366036 661194
rect 6269 661136 6274 661192
rect 6330 661136 366036 661192
rect 6269 661134 366036 661136
rect 6269 661131 6335 661134
rect 366030 661132 366036 661134
rect 366100 661132 366106 661196
rect 98678 660996 98684 661060
rect 98748 661058 98754 661060
rect 545614 661058 545620 661060
rect 98748 660998 545620 661058
rect 98748 660996 98754 660998
rect 545614 660996 545620 660998
rect 545684 660996 545690 661060
rect 53598 660860 53604 660924
rect 53668 660922 53674 660924
rect 66294 660922 66300 660924
rect 53668 660862 66300 660922
rect 53668 660860 53674 660862
rect 66294 660860 66300 660862
rect 66364 660860 66370 660924
rect 333830 660860 333836 660924
rect 333900 660922 333906 660924
rect 352046 660922 352052 660924
rect 333900 660862 352052 660922
rect 333900 660860 333906 660862
rect 352046 660860 352052 660862
rect 352116 660860 352122 660924
rect 542077 660922 542143 660925
rect 544326 660922 544332 660924
rect 542077 660920 544332 660922
rect 542077 660864 542082 660920
rect 542138 660864 544332 660920
rect 542077 660862 544332 660864
rect 542077 660859 542143 660862
rect 544326 660860 544332 660862
rect 544396 660860 544402 660924
rect 35157 660786 35223 660789
rect 108982 660786 108988 660788
rect 35157 660784 108988 660786
rect 35157 660728 35162 660784
rect 35218 660728 108988 660784
rect 35157 660726 108988 660728
rect 35157 660723 35223 660726
rect 108982 660724 108988 660726
rect 109052 660724 109058 660788
rect 310462 660724 310468 660788
rect 310532 660786 310538 660788
rect 352230 660786 352236 660788
rect 310532 660726 352236 660786
rect 310532 660724 310538 660726
rect 352230 660724 352236 660726
rect 352300 660724 352306 660788
rect 39389 660650 39455 660653
rect 121494 660650 121500 660652
rect 39389 660648 121500 660650
rect 39389 660592 39394 660648
rect 39450 660592 121500 660648
rect 39389 660590 121500 660592
rect 39389 660587 39455 660590
rect 121494 660588 121500 660590
rect 121564 660588 121570 660652
rect 301446 660588 301452 660652
rect 301516 660650 301522 660652
rect 353518 660650 353524 660652
rect 301516 660590 353524 660650
rect 301516 660588 301522 660590
rect 353518 660588 353524 660590
rect 353588 660588 353594 660652
rect 40953 660514 41019 660517
rect 46238 660514 46244 660516
rect 40953 660512 46244 660514
rect 40953 660456 40958 660512
rect 41014 660456 46244 660512
rect 40953 660454 46244 660456
rect 40953 660451 41019 660454
rect 46238 660452 46244 660454
rect 46308 660452 46314 660516
rect 54702 660452 54708 660516
rect 54772 660514 54778 660516
rect 172462 660514 172468 660516
rect 54772 660454 172468 660514
rect 54772 660452 54778 660454
rect 172462 660452 172468 660454
rect 172532 660452 172538 660516
rect 285806 660452 285812 660516
rect 285876 660514 285882 660516
rect 352414 660514 352420 660516
rect 285876 660454 352420 660514
rect 285876 660452 285882 660454
rect 352414 660452 352420 660454
rect 352484 660452 352490 660516
rect 542537 660514 542603 660517
rect 543590 660514 543596 660516
rect 542537 660512 543596 660514
rect 542537 660456 542542 660512
rect 542598 660456 543596 660512
rect 542537 660454 543596 660456
rect 542537 660451 542603 660454
rect 543590 660452 543596 660454
rect 543660 660452 543666 660516
rect 41505 660378 41571 660381
rect 49734 660378 49740 660380
rect 41505 660376 49740 660378
rect 41505 660320 41510 660376
rect 41566 660320 49740 660376
rect 41505 660318 49740 660320
rect 41505 660315 41571 660318
rect 49734 660316 49740 660318
rect 49804 660316 49810 660380
rect 54886 660316 54892 660380
rect 54956 660378 54962 660380
rect 179454 660378 179460 660380
rect 54956 660318 179460 660378
rect 54956 660316 54962 660318
rect 179454 660316 179460 660318
rect 179524 660316 179530 660380
rect 297950 660316 297956 660380
rect 298020 660378 298026 660380
rect 425094 660378 425100 660380
rect 298020 660318 425100 660378
rect 298020 660316 298026 660318
rect 425094 660316 425100 660318
rect 425164 660316 425170 660380
rect 544510 660378 544516 660380
rect 528510 660318 544516 660378
rect 10961 660242 11027 660245
rect 528510 660242 528570 660318
rect 544510 660316 544516 660318
rect 544580 660316 544586 660380
rect 10961 660240 528570 660242
rect 10961 660184 10966 660240
rect 11022 660184 528570 660240
rect 10961 660182 528570 660184
rect 10961 660179 11027 660182
rect 542118 660180 542124 660244
rect 542188 660180 542194 660244
rect 542302 660180 542308 660244
rect 542372 660180 542378 660244
rect 41689 660106 41755 660109
rect 542126 660106 542186 660180
rect 41689 660104 542186 660106
rect 41689 660048 41694 660104
rect 41750 660048 542186 660104
rect 41689 660046 542186 660048
rect 41689 660043 41755 660046
rect 46238 659908 46244 659972
rect 46308 659970 46314 659972
rect 542310 659970 542370 660180
rect 46308 659910 542370 659970
rect 46308 659908 46314 659910
rect 38745 659834 38811 659837
rect 38745 659832 41124 659834
rect 38745 659776 38750 659832
rect 38806 659776 41124 659832
rect 38745 659774 41124 659776
rect 38745 659771 38811 659774
rect 544653 659562 544719 659565
rect 542892 659560 544719 659562
rect -960 659426 480 659516
rect 542892 659504 544658 659560
rect 544714 659504 544719 659560
rect 542892 659502 544719 659504
rect 544653 659499 544719 659502
rect 3417 659426 3483 659429
rect -960 659424 3483 659426
rect -960 659368 3422 659424
rect 3478 659368 3483 659424
rect -960 659366 3483 659368
rect -960 659276 480 659366
rect 3417 659363 3483 659366
rect 39297 657388 39363 657389
rect 39246 657386 39252 657388
rect 39206 657326 39252 657386
rect 39316 657384 39363 657388
rect 39358 657328 39363 657384
rect 39246 657324 39252 657326
rect 39316 657324 39363 657328
rect 39297 657323 39363 657324
rect 580809 657250 580875 657253
rect 583520 657250 584960 657340
rect 580809 657248 584960 657250
rect 580809 657192 580814 657248
rect 580870 657192 584960 657248
rect 580809 657190 584960 657192
rect 580809 657187 580875 657190
rect 583520 657100 584960 657190
rect 38837 655482 38903 655485
rect 38837 655480 41124 655482
rect 38837 655424 38842 655480
rect 38898 655424 41124 655480
rect 38837 655422 41124 655424
rect 38837 655419 38903 655422
rect 544009 655210 544075 655213
rect 542892 655208 544075 655210
rect 542892 655152 544014 655208
rect 544070 655152 544075 655208
rect 542892 655150 544075 655152
rect 544009 655147 544075 655150
rect -960 654530 480 654620
rect 3417 654530 3483 654533
rect -960 654528 3483 654530
rect -960 654472 3422 654528
rect 3478 654472 3483 654528
rect -960 654470 3483 654472
rect -960 654380 480 654470
rect 3417 654467 3483 654470
rect 542118 653380 542124 653444
rect 542188 653442 542194 653444
rect 562317 653442 562383 653445
rect 542188 653440 562383 653442
rect 542188 653384 562322 653440
rect 562378 653384 562383 653440
rect 542188 653382 562383 653384
rect 542188 653380 542194 653382
rect 562317 653379 562383 653382
rect 580625 652354 580691 652357
rect 583520 652354 584960 652444
rect 580625 652352 584960 652354
rect 580625 652296 580630 652352
rect 580686 652296 584960 652352
rect 580625 652294 584960 652296
rect 580625 652291 580691 652294
rect 583520 652204 584960 652294
rect 543641 651130 543707 651133
rect 542862 651128 543707 651130
rect 542862 651072 543646 651128
rect 543702 651072 543707 651128
rect 542862 651070 543707 651072
rect 38837 650858 38903 650861
rect 38837 650856 41124 650858
rect 38837 650800 38842 650856
rect 38898 650800 41124 650856
rect 38837 650798 41124 650800
rect 38837 650795 38903 650798
rect 542862 650556 542922 651070
rect 543641 651067 543707 651070
rect -960 649634 480 649724
rect 3325 649634 3391 649637
rect -960 649632 3391 649634
rect -960 649576 3330 649632
rect 3386 649576 3391 649632
rect -960 649574 3391 649576
rect -960 649484 480 649574
rect 3325 649571 3391 649574
rect 583520 647036 584960 647276
rect 38837 646506 38903 646509
rect 38837 646504 41124 646506
rect 38837 646448 38842 646504
rect 38898 646448 41124 646504
rect 38837 646446 41124 646448
rect 38837 646443 38903 646446
rect 544837 646234 544903 646237
rect 542892 646232 544903 646234
rect 542892 646176 544842 646232
rect 544898 646176 544903 646232
rect 542892 646174 544903 646176
rect 544837 646171 544903 646174
rect -960 644466 480 644556
rect 3693 644466 3759 644469
rect -960 644464 3759 644466
rect -960 644408 3698 644464
rect 3754 644408 3759 644464
rect -960 644406 3759 644408
rect -960 644316 480 644406
rect 3693 644403 3759 644406
rect 580073 642290 580139 642293
rect 583520 642290 584960 642380
rect 580073 642288 584960 642290
rect 580073 642232 580078 642288
rect 580134 642232 584960 642288
rect 580073 642230 584960 642232
rect 580073 642227 580139 642230
rect 583520 642140 584960 642230
rect 38837 641882 38903 641885
rect 542721 641882 542787 641885
rect 38837 641880 41124 641882
rect 38837 641824 38842 641880
rect 38898 641824 41124 641880
rect 38837 641822 41124 641824
rect 542678 641880 542787 641882
rect 542678 641824 542726 641880
rect 542782 641824 542787 641880
rect 38837 641819 38903 641822
rect 542678 641819 542787 641824
rect 542678 641580 542738 641819
rect -960 639570 480 639660
rect 2773 639570 2839 639573
rect -960 639568 2839 639570
rect -960 639512 2778 639568
rect 2834 639512 2839 639568
rect -960 639510 2839 639512
rect -960 639420 480 639510
rect 2773 639507 2839 639510
rect 39757 637530 39823 637533
rect 39757 637528 41124 637530
rect 39757 637472 39762 637528
rect 39818 637472 41124 637528
rect 39757 637470 41124 637472
rect 39757 637467 39823 637470
rect 579981 637394 580047 637397
rect 583520 637394 584960 637484
rect 579981 637392 584960 637394
rect 579981 637336 579986 637392
rect 580042 637336 584960 637392
rect 579981 637334 584960 637336
rect 579981 637331 580047 637334
rect 544837 637258 544903 637261
rect 542892 637256 544903 637258
rect 542892 637200 544842 637256
rect 544898 637200 544903 637256
rect 583520 637244 584960 637334
rect 542892 637198 544903 637200
rect 544837 637195 544903 637198
rect -960 634674 480 634764
rect 2773 634674 2839 634677
rect -960 634672 2839 634674
rect -960 634616 2778 634672
rect 2834 634616 2839 634672
rect -960 634614 2839 634616
rect -960 634524 480 634614
rect 2773 634611 2839 634614
rect 542629 633450 542695 633453
rect 542629 633448 542738 633450
rect 542629 633392 542634 633448
rect 542690 633392 542738 633448
rect 542629 633387 542738 633392
rect 39941 632906 40007 632909
rect 39941 632904 41124 632906
rect 39941 632848 39946 632904
rect 40002 632848 41124 632904
rect 542678 632876 542738 633387
rect 39941 632846 41124 632848
rect 39941 632843 40007 632846
rect 580165 632498 580231 632501
rect 583520 632498 584960 632588
rect 580165 632496 584960 632498
rect 580165 632440 580170 632496
rect 580226 632440 584960 632496
rect 580165 632438 584960 632440
rect 580165 632435 580231 632438
rect 583520 632348 584960 632438
rect -960 629778 480 629868
rect 3509 629778 3575 629781
rect -960 629776 3575 629778
rect -960 629720 3514 629776
rect 3570 629720 3575 629776
rect -960 629718 3575 629720
rect -960 629628 480 629718
rect 3509 629715 3575 629718
rect 38929 628418 38995 628421
rect 38929 628416 41124 628418
rect 38929 628360 38934 628416
rect 38990 628360 41124 628416
rect 38929 628358 41124 628360
rect 38929 628355 38995 628358
rect 544101 628146 544167 628149
rect 542892 628144 544167 628146
rect 542892 628088 544106 628144
rect 544162 628088 544167 628144
rect 542892 628086 544167 628088
rect 544101 628083 544167 628086
rect 583520 627452 584960 627692
rect -960 624882 480 624972
rect 3877 624882 3943 624885
rect -960 624880 3943 624882
rect -960 624824 3882 624880
rect 3938 624824 3943 624880
rect -960 624822 3943 624824
rect -960 624732 480 624822
rect 3877 624819 3943 624822
rect 544837 623930 544903 623933
rect 542892 623928 544903 623930
rect 542892 623872 544842 623928
rect 544898 623872 544903 623928
rect 542892 623870 544903 623872
rect 544837 623867 544903 623870
rect 39798 623732 39804 623796
rect 39868 623794 39874 623796
rect 39868 623734 41124 623794
rect 39868 623732 39874 623734
rect 580165 622706 580231 622709
rect 583520 622706 584960 622796
rect 580165 622704 584960 622706
rect 580165 622648 580170 622704
rect 580226 622648 584960 622704
rect 580165 622646 584960 622648
rect 580165 622643 580231 622646
rect 583520 622556 584960 622646
rect -960 619836 480 620076
rect 38837 619442 38903 619445
rect 38837 619440 41124 619442
rect 38837 619384 38842 619440
rect 38898 619384 41124 619440
rect 38837 619382 41124 619384
rect 38837 619379 38903 619382
rect 544837 619170 544903 619173
rect 542892 619168 544903 619170
rect 542892 619112 544842 619168
rect 544898 619112 544903 619168
rect 542892 619110 544903 619112
rect 544837 619107 544903 619110
rect 579981 617810 580047 617813
rect 583520 617810 584960 617900
rect 579981 617808 584960 617810
rect 579981 617752 579986 617808
rect 580042 617752 584960 617808
rect 579981 617750 584960 617752
rect 579981 617747 580047 617750
rect 583520 617660 584960 617750
rect 542629 615226 542695 615229
rect 542629 615224 542738 615226
rect -960 615090 480 615180
rect 542629 615168 542634 615224
rect 542690 615168 542738 615224
rect 542629 615163 542738 615168
rect 3325 615090 3391 615093
rect -960 615088 3391 615090
rect -960 615032 3330 615088
rect 3386 615032 3391 615088
rect -960 615030 3391 615032
rect -960 614940 480 615030
rect 3325 615027 3391 615030
rect 38837 615090 38903 615093
rect 38837 615088 41124 615090
rect 38837 615032 38842 615088
rect 38898 615032 41124 615088
rect 38837 615030 41124 615032
rect 38837 615027 38903 615030
rect 542678 614924 542738 615163
rect 579613 612914 579679 612917
rect 583520 612914 584960 613004
rect 579613 612912 584960 612914
rect 579613 612856 579618 612912
rect 579674 612856 584960 612912
rect 579613 612854 584960 612856
rect 579613 612851 579679 612854
rect 583520 612764 584960 612854
rect 541985 610874 542051 610877
rect 541942 610872 542051 610874
rect 541942 610816 541990 610872
rect 542046 610816 542051 610872
rect 541942 610811 542051 610816
rect 39430 610404 39436 610468
rect 39500 610466 39506 610468
rect 39500 610406 41124 610466
rect 39500 610404 39506 610406
rect 541942 610300 542002 610811
rect -960 610194 480 610284
rect 3325 610194 3391 610197
rect -960 610192 3391 610194
rect -960 610136 3330 610192
rect 3386 610136 3391 610192
rect -960 610134 3391 610136
rect -960 610044 480 610134
rect 3325 610131 3391 610134
rect 580165 608018 580231 608021
rect 583520 608018 584960 608108
rect 580165 608016 584960 608018
rect 580165 607960 580170 608016
rect 580226 607960 584960 608016
rect 580165 607958 584960 607960
rect 580165 607955 580231 607958
rect 583520 607868 584960 607958
rect 39246 606188 39252 606252
rect 39316 606250 39322 606252
rect 39316 606190 41124 606250
rect 39316 606188 39322 606190
rect 544837 605978 544903 605981
rect 542892 605976 544903 605978
rect 542892 605920 544842 605976
rect 544898 605920 544903 605976
rect 542892 605918 544903 605920
rect 544837 605915 544903 605918
rect -960 605298 480 605388
rect 3325 605298 3391 605301
rect -960 605296 3391 605298
rect -960 605240 3330 605296
rect 3386 605240 3391 605296
rect -960 605238 3391 605240
rect -960 605148 480 605238
rect 3325 605235 3391 605238
rect 579613 603122 579679 603125
rect 583520 603122 584960 603212
rect 579613 603120 584960 603122
rect 579613 603064 579618 603120
rect 579674 603064 584960 603120
rect 579613 603062 584960 603064
rect 579613 603059 579679 603062
rect 583520 602972 584960 603062
rect 38837 601626 38903 601629
rect 38837 601624 41124 601626
rect 38837 601568 38842 601624
rect 38898 601568 41124 601624
rect 38837 601566 41124 601568
rect 38837 601563 38903 601566
rect 544837 601218 544903 601221
rect 542892 601216 544903 601218
rect 542892 601160 544842 601216
rect 544898 601160 544903 601216
rect 542892 601158 544903 601160
rect 544837 601155 544903 601158
rect -960 600402 480 600492
rect 2773 600402 2839 600405
rect -960 600400 2839 600402
rect -960 600344 2778 600400
rect 2834 600344 2839 600400
rect -960 600342 2839 600344
rect -960 600252 480 600342
rect 2773 600339 2839 600342
rect 580165 598226 580231 598229
rect 583520 598226 584960 598316
rect 580165 598224 584960 598226
rect 580165 598168 580170 598224
rect 580226 598168 584960 598224
rect 580165 598166 584960 598168
rect 580165 598163 580231 598166
rect 583520 598076 584960 598166
rect 38837 597274 38903 597277
rect 38837 597272 41124 597274
rect 38837 597216 38842 597272
rect 38898 597216 41124 597272
rect 38837 597214 41124 597216
rect 38837 597211 38903 597214
rect 543641 597002 543707 597005
rect 542892 597000 543707 597002
rect 542892 596944 543646 597000
rect 543702 596944 543707 597000
rect 542892 596942 543707 596944
rect 543641 596939 543707 596942
rect -960 595506 480 595596
rect 3325 595506 3391 595509
rect -960 595504 3391 595506
rect -960 595448 3330 595504
rect 3386 595448 3391 595504
rect -960 595446 3391 595448
rect -960 595356 480 595446
rect 3325 595443 3391 595446
rect 579613 593058 579679 593061
rect 583520 593058 584960 593148
rect 579613 593056 584960 593058
rect 579613 593000 579618 593056
rect 579674 593000 584960 593056
rect 579613 592998 584960 593000
rect 579613 592995 579679 592998
rect 542302 592860 542308 592924
rect 542372 592860 542378 592924
rect 583520 592908 584960 592998
rect 38837 592514 38903 592517
rect 38837 592512 41124 592514
rect 38837 592456 38842 592512
rect 38898 592456 41124 592512
rect 38837 592454 41124 592456
rect 38837 592451 38903 592454
rect 542310 592348 542370 592860
rect -960 590338 480 590428
rect 3141 590338 3207 590341
rect -960 590336 3207 590338
rect -960 590280 3146 590336
rect 3202 590280 3207 590336
rect -960 590278 3207 590280
rect -960 590188 480 590278
rect 3141 590275 3207 590278
rect 38837 588298 38903 588301
rect 38837 588296 41124 588298
rect 38837 588240 38842 588296
rect 38898 588240 41124 588296
rect 38837 588238 41124 588240
rect 38837 588235 38903 588238
rect 580165 588162 580231 588165
rect 583520 588162 584960 588252
rect 580165 588160 584960 588162
rect 580165 588104 580170 588160
rect 580226 588104 584960 588160
rect 580165 588102 584960 588104
rect 580165 588099 580231 588102
rect 583520 588012 584960 588102
rect 542310 587756 542370 587860
rect 542302 587692 542308 587756
rect 542372 587692 542378 587756
rect -960 585442 480 585532
rect 2773 585442 2839 585445
rect -960 585440 2839 585442
rect -960 585384 2778 585440
rect 2834 585384 2839 585440
rect -960 585382 2839 585384
rect -960 585292 480 585382
rect 2773 585379 2839 585382
rect 40125 583674 40191 583677
rect 40125 583672 41124 583674
rect 40125 583616 40130 583672
rect 40186 583616 41124 583672
rect 40125 583614 41124 583616
rect 40125 583611 40191 583614
rect 545246 583266 545252 583268
rect 542892 583206 545252 583266
rect 545246 583204 545252 583206
rect 545316 583204 545322 583268
rect 579981 583266 580047 583269
rect 583520 583266 584960 583356
rect 579981 583264 584960 583266
rect 579981 583208 579986 583264
rect 580042 583208 584960 583264
rect 579981 583206 584960 583208
rect 579981 583203 580047 583206
rect 583520 583116 584960 583206
rect 39757 582450 39823 582453
rect 40534 582450 40540 582452
rect 39757 582448 40540 582450
rect 39757 582392 39762 582448
rect 39818 582392 40540 582448
rect 39757 582390 40540 582392
rect 39757 582387 39823 582390
rect 40534 582388 40540 582390
rect 40604 582388 40610 582452
rect -960 580546 480 580636
rect 3233 580546 3299 580549
rect -960 580544 3299 580546
rect -960 580488 3238 580544
rect 3294 580488 3299 580544
rect -960 580486 3299 580488
rect -960 580396 480 580486
rect 3233 580483 3299 580486
rect 39021 579322 39087 579325
rect 39021 579320 41124 579322
rect 39021 579264 39026 579320
rect 39082 579264 41124 579320
rect 39021 579262 41124 579264
rect 39021 579259 39087 579262
rect 542862 578370 542922 578884
rect 545297 578370 545363 578373
rect 542862 578368 545363 578370
rect 542862 578312 545302 578368
rect 545358 578312 545363 578368
rect 542862 578310 545363 578312
rect 545297 578307 545363 578310
rect 579613 578370 579679 578373
rect 583520 578370 584960 578460
rect 579613 578368 584960 578370
rect 579613 578312 579618 578368
rect 579674 578312 584960 578368
rect 579613 578310 584960 578312
rect 579613 578307 579679 578310
rect 583520 578220 584960 578310
rect -960 575650 480 575740
rect 3141 575650 3207 575653
rect -960 575648 3207 575650
rect -960 575592 3146 575648
rect 3202 575592 3207 575648
rect -960 575590 3207 575592
rect -960 575500 480 575590
rect 3141 575587 3207 575590
rect 544929 574698 544995 574701
rect 542892 574696 544995 574698
rect 542892 574640 544934 574696
rect 544990 574640 544995 574696
rect 542892 574638 544995 574640
rect 544929 574635 544995 574638
rect 38837 574562 38903 574565
rect 38837 574560 41124 574562
rect 38837 574504 38842 574560
rect 38898 574504 41124 574560
rect 38837 574502 41124 574504
rect 38837 574499 38903 574502
rect 580165 573474 580231 573477
rect 583520 573474 584960 573564
rect 580165 573472 584960 573474
rect 580165 573416 580170 573472
rect 580226 573416 584960 573472
rect 580165 573414 584960 573416
rect 580165 573411 580231 573414
rect 583520 573324 584960 573414
rect -960 570754 480 570844
rect 3049 570754 3115 570757
rect -960 570752 3115 570754
rect -960 570696 3054 570752
rect 3110 570696 3115 570752
rect -960 570694 3115 570696
rect -960 570604 480 570694
rect 3049 570691 3115 570694
rect 39113 570346 39179 570349
rect 39113 570344 41124 570346
rect 39113 570288 39118 570344
rect 39174 570288 41124 570344
rect 39113 570286 41124 570288
rect 39113 570283 39179 570286
rect 544929 570074 544995 570077
rect 542892 570072 544995 570074
rect 542892 570016 544934 570072
rect 544990 570016 544995 570072
rect 542892 570014 544995 570016
rect 544929 570011 544995 570014
rect 583520 568428 584960 568668
rect -960 565858 480 565948
rect 2773 565858 2839 565861
rect -960 565856 2839 565858
rect -960 565800 2778 565856
rect 2834 565800 2839 565856
rect -960 565798 2839 565800
rect -960 565708 480 565798
rect 2773 565795 2839 565798
rect 38653 565722 38719 565725
rect 544929 565722 544995 565725
rect 38653 565720 41124 565722
rect 38653 565664 38658 565720
rect 38714 565664 41124 565720
rect 38653 565662 41124 565664
rect 542892 565720 544995 565722
rect 542892 565664 544934 565720
rect 544990 565664 544995 565720
rect 542892 565662 544995 565664
rect 38653 565659 38719 565662
rect 544929 565659 544995 565662
rect 583520 563532 584960 563772
rect 38653 561370 38719 561373
rect 38653 561368 41124 561370
rect 38653 561312 38658 561368
rect 38714 561312 41124 561368
rect 38653 561310 41124 561312
rect 38653 561307 38719 561310
rect 545021 561098 545087 561101
rect 542892 561096 545087 561098
rect -960 560962 480 561052
rect 542892 561040 545026 561096
rect 545082 561040 545087 561096
rect 542892 561038 545087 561040
rect 545021 561035 545087 561038
rect 3141 560962 3207 560965
rect -960 560960 3207 560962
rect -960 560904 3146 560960
rect 3202 560904 3207 560960
rect -960 560902 3207 560904
rect -960 560812 480 560902
rect 3141 560899 3207 560902
rect 580165 558786 580231 558789
rect 583520 558786 584960 558876
rect 580165 558784 584960 558786
rect 580165 558728 580170 558784
rect 580226 558728 584960 558784
rect 580165 558726 584960 558728
rect 580165 558723 580231 558726
rect 583520 558636 584960 558726
rect 38653 556882 38719 556885
rect 38653 556880 41124 556882
rect 38653 556824 38658 556880
rect 38714 556824 41124 556880
rect 38653 556822 41124 556824
rect 38653 556819 38719 556822
rect 545297 556610 545363 556613
rect 542892 556608 545363 556610
rect 542892 556552 545302 556608
rect 545358 556552 545363 556608
rect 542892 556550 545363 556552
rect 545297 556547 545363 556550
rect -960 556066 480 556156
rect 3141 556066 3207 556069
rect -960 556064 3207 556066
rect -960 556008 3146 556064
rect 3202 556008 3207 556064
rect -960 556006 3207 556008
rect -960 555916 480 556006
rect 3141 556003 3207 556006
rect 580165 553890 580231 553893
rect 583520 553890 584960 553980
rect 580165 553888 584960 553890
rect 580165 553832 580170 553888
rect 580226 553832 584960 553888
rect 580165 553830 584960 553832
rect 580165 553827 580231 553830
rect 583520 553740 584960 553830
rect 39941 552394 40007 552397
rect 39941 552392 41124 552394
rect 39941 552336 39946 552392
rect 40002 552336 41124 552392
rect 39941 552334 41124 552336
rect 39941 552331 40007 552334
rect 544929 552122 544995 552125
rect 542892 552120 544995 552122
rect 542892 552064 544934 552120
rect 544990 552064 544995 552120
rect 542892 552062 544995 552064
rect 544929 552059 544995 552062
rect -960 551170 480 551260
rect 3141 551170 3207 551173
rect -960 551168 3207 551170
rect -960 551112 3146 551168
rect 3202 551112 3207 551168
rect -960 551110 3207 551112
rect -960 551020 480 551110
rect 3141 551107 3207 551110
rect 580533 548994 580599 548997
rect 583520 548994 584960 549084
rect 580533 548992 584960 548994
rect 580533 548936 580538 548992
rect 580594 548936 584960 548992
rect 580533 548934 584960 548936
rect 580533 548931 580599 548934
rect 583520 548844 584960 548934
rect 39205 548042 39271 548045
rect 39205 548040 41124 548042
rect 39205 547984 39210 548040
rect 39266 547984 41124 548040
rect 39205 547982 41124 547984
rect 39205 547979 39271 547982
rect 544653 547634 544719 547637
rect 542892 547632 544719 547634
rect 542892 547576 544658 547632
rect 544714 547576 544719 547632
rect 542892 547574 544719 547576
rect 544653 547571 544719 547574
rect -960 546274 480 546364
rect 3141 546274 3207 546277
rect -960 546272 3207 546274
rect -960 546216 3146 546272
rect 3202 546216 3207 546272
rect -960 546214 3207 546216
rect -960 546124 480 546214
rect 3141 546211 3207 546214
rect 580073 544098 580139 544101
rect 583520 544098 584960 544188
rect 580073 544096 584960 544098
rect 580073 544040 580078 544096
rect 580134 544040 584960 544096
rect 580073 544038 584960 544040
rect 580073 544035 580139 544038
rect 583520 543948 584960 544038
rect 38009 543418 38075 543421
rect 38009 543416 41124 543418
rect 38009 543360 38014 543416
rect 38070 543360 41124 543416
rect 38009 543358 41124 543360
rect 38009 543355 38075 543358
rect 543958 543010 543964 543012
rect 542892 542950 543964 543010
rect 543958 542948 543964 542950
rect 544028 542948 544034 543012
rect -960 541378 480 541468
rect 3141 541378 3207 541381
rect -960 541376 3207 541378
rect -960 541320 3146 541376
rect 3202 541320 3207 541376
rect -960 541318 3207 541320
rect -960 541228 480 541318
rect 3141 541315 3207 541318
rect 38653 539066 38719 539069
rect 38653 539064 41124 539066
rect 38653 539008 38658 539064
rect 38714 539008 41124 539064
rect 38653 539006 41124 539008
rect 38653 539003 38719 539006
rect 580165 538930 580231 538933
rect 583520 538930 584960 539020
rect 580165 538928 584960 538930
rect 580165 538872 580170 538928
rect 580226 538872 584960 538928
rect 580165 538870 584960 538872
rect 580165 538867 580231 538870
rect 544929 538794 544995 538797
rect 542892 538792 544995 538794
rect 542892 538736 544934 538792
rect 544990 538736 544995 538792
rect 583520 538780 584960 538870
rect 542892 538734 544995 538736
rect 544929 538731 544995 538734
rect -960 536060 480 536300
rect 39941 534442 40007 534445
rect 39941 534440 41124 534442
rect 39941 534384 39946 534440
rect 40002 534384 41124 534440
rect 39941 534382 41124 534384
rect 39941 534379 40007 534382
rect 544653 534170 544719 534173
rect 542892 534168 544719 534170
rect 542892 534112 544658 534168
rect 544714 534112 544719 534168
rect 542892 534110 544719 534112
rect 544653 534107 544719 534110
rect 580257 534034 580323 534037
rect 583520 534034 584960 534124
rect 580257 534032 584960 534034
rect 580257 533976 580262 534032
rect 580318 533976 584960 534032
rect 580257 533974 584960 533976
rect 580257 533971 580323 533974
rect 583520 533884 584960 533974
rect -960 531314 480 531404
rect 2773 531314 2839 531317
rect -960 531312 2839 531314
rect -960 531256 2778 531312
rect 2834 531256 2839 531312
rect -960 531254 2839 531256
rect -960 531164 480 531254
rect 2773 531251 2839 531254
rect 542537 530090 542603 530093
rect 542494 530088 542603 530090
rect 542494 530032 542542 530088
rect 542598 530032 542603 530088
rect 542494 530027 542603 530032
rect 38653 529954 38719 529957
rect 38653 529952 41124 529954
rect 38653 529896 38658 529952
rect 38714 529896 41124 529952
rect 38653 529894 41124 529896
rect 38653 529891 38719 529894
rect 542494 529788 542554 530027
rect 580165 529138 580231 529141
rect 583520 529138 584960 529228
rect 580165 529136 584960 529138
rect 580165 529080 580170 529136
rect 580226 529080 584960 529136
rect 580165 529078 584960 529080
rect 580165 529075 580231 529078
rect 583520 528988 584960 529078
rect -960 526268 480 526508
rect 38653 525466 38719 525469
rect 38653 525464 41124 525466
rect 38653 525408 38658 525464
rect 38714 525408 41124 525464
rect 38653 525406 41124 525408
rect 38653 525403 38719 525406
rect 542494 524517 542554 525028
rect 542494 524512 542603 524517
rect 542494 524456 542542 524512
rect 542598 524456 542603 524512
rect 542494 524454 542603 524456
rect 542537 524451 542603 524454
rect 579613 524242 579679 524245
rect 583520 524242 584960 524332
rect 579613 524240 584960 524242
rect 579613 524184 579618 524240
rect 579674 524184 584960 524240
rect 579613 524182 584960 524184
rect 579613 524179 579679 524182
rect 583520 524092 584960 524182
rect -960 521522 480 521612
rect 3141 521522 3207 521525
rect -960 521520 3207 521522
rect -960 521464 3146 521520
rect 3202 521464 3207 521520
rect -960 521462 3207 521464
rect -960 521372 480 521462
rect 3141 521459 3207 521462
rect 38009 520978 38075 520981
rect 38009 520976 41124 520978
rect 38009 520920 38014 520976
rect 38070 520920 41124 520976
rect 38009 520918 41124 520920
rect 38009 520915 38075 520918
rect 544653 520842 544719 520845
rect 542892 520840 544719 520842
rect 542892 520784 544658 520840
rect 544714 520784 544719 520840
rect 542892 520782 544719 520784
rect 544653 520779 544719 520782
rect 580257 519346 580323 519349
rect 583520 519346 584960 519436
rect 580257 519344 584960 519346
rect 580257 519288 580262 519344
rect 580318 519288 584960 519344
rect 580257 519286 584960 519288
rect 580257 519283 580323 519286
rect 583520 519196 584960 519286
rect -960 516626 480 516716
rect 3693 516626 3759 516629
rect -960 516624 3759 516626
rect -960 516568 3698 516624
rect 3754 516568 3759 516624
rect -960 516566 3759 516568
rect -960 516476 480 516566
rect 3693 516563 3759 516566
rect 39246 516292 39252 516356
rect 39316 516354 39322 516356
rect 545021 516354 545087 516357
rect 39316 516294 41124 516354
rect 542892 516352 545087 516354
rect 542892 516296 545026 516352
rect 545082 516296 545087 516352
rect 542892 516294 545087 516296
rect 39316 516292 39322 516294
rect 545021 516291 545087 516294
rect 580165 514450 580231 514453
rect 583520 514450 584960 514540
rect 580165 514448 584960 514450
rect 580165 514392 580170 514448
rect 580226 514392 584960 514448
rect 580165 514390 584960 514392
rect 580165 514387 580231 514390
rect 583520 514300 584960 514390
rect 38653 512138 38719 512141
rect 38653 512136 41124 512138
rect 38653 512080 38658 512136
rect 38714 512080 41124 512136
rect 38653 512078 41124 512080
rect 38653 512075 38719 512078
rect 544653 511866 544719 511869
rect 542892 511864 544719 511866
rect -960 511730 480 511820
rect 542892 511808 544658 511864
rect 544714 511808 544719 511864
rect 542892 511806 544719 511808
rect 544653 511803 544719 511806
rect 3141 511730 3207 511733
rect -960 511728 3207 511730
rect -960 511672 3146 511728
rect 3202 511672 3207 511728
rect -960 511670 3207 511672
rect -960 511580 480 511670
rect 3141 511667 3207 511670
rect 580533 509554 580599 509557
rect 583520 509554 584960 509644
rect 580533 509552 584960 509554
rect 580533 509496 580538 509552
rect 580594 509496 584960 509552
rect 580533 509494 584960 509496
rect 580533 509491 580599 509494
rect 583520 509404 584960 509494
rect 40125 507378 40191 507381
rect 544653 507378 544719 507381
rect 40125 507376 41124 507378
rect 40125 507320 40130 507376
rect 40186 507320 41124 507376
rect 40125 507318 41124 507320
rect 542892 507376 544719 507378
rect 542892 507320 544658 507376
rect 544714 507320 544719 507376
rect 542892 507318 544719 507320
rect 40125 507315 40191 507318
rect 544653 507315 544719 507318
rect -960 506834 480 506924
rect 3509 506834 3575 506837
rect -960 506832 3575 506834
rect -960 506776 3514 506832
rect 3570 506776 3575 506832
rect -960 506774 3575 506776
rect -960 506684 480 506774
rect 3509 506771 3575 506774
rect 579981 504658 580047 504661
rect 583520 504658 584960 504748
rect 579981 504656 584960 504658
rect 579981 504600 579986 504656
rect 580042 504600 584960 504656
rect 579981 504598 584960 504600
rect 579981 504595 580047 504598
rect 583520 504508 584960 504598
rect 542629 503434 542695 503437
rect 542629 503432 542738 503434
rect 542629 503376 542634 503432
rect 542690 503376 542738 503432
rect 542629 503371 542738 503376
rect 38745 503162 38811 503165
rect 38745 503160 41124 503162
rect 38745 503104 38750 503160
rect 38806 503104 41124 503160
rect 38745 503102 41124 503104
rect 38745 503099 38811 503102
rect 542678 502860 542738 503371
rect -960 501938 480 502028
rect 3693 501938 3759 501941
rect -960 501936 3759 501938
rect -960 501880 3698 501936
rect 3754 501880 3759 501936
rect -960 501878 3759 501880
rect -960 501788 480 501878
rect 3693 501875 3759 501878
rect 579705 499762 579771 499765
rect 583520 499762 584960 499852
rect 579705 499760 584960 499762
rect 579705 499704 579710 499760
rect 579766 499704 584960 499760
rect 579705 499702 584960 499704
rect 579705 499699 579771 499702
rect 583520 499612 584960 499702
rect 38745 498810 38811 498813
rect 38745 498808 41124 498810
rect 38745 498752 38750 498808
rect 38806 498752 41124 498808
rect 38745 498750 41124 498752
rect 38745 498747 38811 498750
rect 545021 498402 545087 498405
rect 542892 498400 545087 498402
rect 542892 498344 545026 498400
rect 545082 498344 545087 498400
rect 542892 498342 545087 498344
rect 545021 498339 545087 498342
rect -960 497042 480 497132
rect 3693 497042 3759 497045
rect -960 497040 3759 497042
rect -960 496984 3698 497040
rect 3754 496984 3759 497040
rect -960 496982 3759 496984
rect -960 496892 480 496982
rect 3693 496979 3759 496982
rect 579981 494866 580047 494869
rect 583520 494866 584960 494956
rect 579981 494864 584960 494866
rect 579981 494808 579986 494864
rect 580042 494808 584960 494864
rect 579981 494806 584960 494808
rect 579981 494803 580047 494806
rect 583520 494716 584960 494806
rect 38745 494186 38811 494189
rect 38745 494184 41124 494186
rect 38745 494128 38750 494184
rect 38806 494128 41124 494184
rect 38745 494126 41124 494128
rect 38745 494123 38811 494126
rect 544653 493914 544719 493917
rect 542892 493912 544719 493914
rect 542892 493856 544658 493912
rect 544714 493856 544719 493912
rect 542892 493854 544719 493856
rect 544653 493851 544719 493854
rect -960 492146 480 492236
rect 3509 492146 3575 492149
rect -960 492144 3575 492146
rect -960 492088 3514 492144
rect 3570 492088 3575 492144
rect -960 492086 3575 492088
rect -960 491996 480 492086
rect 3509 492083 3575 492086
rect 580165 489970 580231 489973
rect 583520 489970 584960 490060
rect 580165 489968 584960 489970
rect 580165 489912 580170 489968
rect 580226 489912 584960 489968
rect 580165 489910 584960 489912
rect 580165 489907 580231 489910
rect 583520 489820 584960 489910
rect 38745 489698 38811 489701
rect 38745 489696 41124 489698
rect 38745 489640 38750 489696
rect 38806 489640 41124 489696
rect 38745 489638 41124 489640
rect 38745 489635 38811 489638
rect 544653 489562 544719 489565
rect 542892 489560 544719 489562
rect 542892 489504 544658 489560
rect 544714 489504 544719 489560
rect 542892 489502 544719 489504
rect 544653 489499 544719 489502
rect -960 487250 480 487340
rect 3141 487250 3207 487253
rect -960 487248 3207 487250
rect -960 487192 3146 487248
rect 3202 487192 3207 487248
rect -960 487190 3207 487192
rect -960 487100 480 487190
rect 3141 487187 3207 487190
rect 38745 485210 38811 485213
rect 38745 485208 41124 485210
rect 38745 485152 38750 485208
rect 38806 485152 41124 485208
rect 38745 485150 41124 485152
rect 38745 485147 38811 485150
rect 580165 484802 580231 484805
rect 583520 484802 584960 484892
rect 580165 484800 584960 484802
rect 542678 484533 542738 484772
rect 580165 484744 580170 484800
rect 580226 484744 584960 484800
rect 580165 484742 584960 484744
rect 580165 484739 580231 484742
rect 583520 484652 584960 484742
rect 542678 484528 542787 484533
rect 542678 484472 542726 484528
rect 542782 484472 542787 484528
rect 542678 484470 542787 484472
rect 542721 484467 542787 484470
rect -960 482082 480 482172
rect 542118 482156 542124 482220
rect 542188 482218 542194 482220
rect 550817 482218 550883 482221
rect 542188 482216 550883 482218
rect 542188 482160 550822 482216
rect 550878 482160 550883 482216
rect 542188 482158 550883 482160
rect 542188 482156 542194 482158
rect 550817 482155 550883 482158
rect 3049 482082 3115 482085
rect -960 482080 3115 482082
rect -960 482024 3054 482080
rect 3110 482024 3115 482080
rect -960 482022 3115 482024
rect -960 481932 480 482022
rect 3049 482019 3115 482022
rect 37917 480722 37983 480725
rect 37917 480720 41124 480722
rect 37917 480664 37922 480720
rect 37978 480664 41124 480720
rect 37917 480662 41124 480664
rect 37917 480659 37983 480662
rect 542678 480317 542738 480420
rect 542629 480312 542738 480317
rect 542629 480256 542634 480312
rect 542690 480256 542738 480312
rect 542629 480254 542738 480256
rect 542629 480251 542695 480254
rect 579613 479906 579679 479909
rect 583520 479906 584960 479996
rect 579613 479904 584960 479906
rect 579613 479848 579618 479904
rect 579674 479848 584960 479904
rect 579613 479846 584960 479848
rect 579613 479843 579679 479846
rect 583520 479756 584960 479846
rect -960 477186 480 477276
rect 2957 477186 3023 477189
rect -960 477184 3023 477186
rect -960 477128 2962 477184
rect 3018 477128 3023 477184
rect -960 477126 3023 477128
rect -960 477036 480 477126
rect 2957 477123 3023 477126
rect 41597 476778 41663 476781
rect 41597 476776 41706 476778
rect 41597 476720 41602 476776
rect 41658 476720 41706 476776
rect 41597 476715 41706 476720
rect 41646 476204 41706 476715
rect 544193 475962 544259 475965
rect 542892 475960 544259 475962
rect 542892 475904 544198 475960
rect 544254 475904 544259 475960
rect 542892 475902 544259 475904
rect 544193 475899 544259 475902
rect 580165 475010 580231 475013
rect 583520 475010 584960 475100
rect 580165 475008 584960 475010
rect 580165 474952 580170 475008
rect 580226 474952 584960 475008
rect 580165 474950 584960 474952
rect 580165 474947 580231 474950
rect 583520 474860 584960 474950
rect -960 472290 480 472380
rect 3509 472290 3575 472293
rect -960 472288 3575 472290
rect -960 472232 3514 472288
rect 3570 472232 3575 472288
rect -960 472230 3575 472232
rect -960 472140 480 472230
rect 3509 472227 3575 472230
rect 39113 471882 39179 471885
rect 541985 471884 542051 471885
rect 39113 471880 41124 471882
rect 39113 471824 39118 471880
rect 39174 471824 41124 471880
rect 39113 471822 41124 471824
rect 39113 471819 39179 471822
rect 541934 471820 541940 471884
rect 542004 471882 542051 471884
rect 542004 471880 542096 471882
rect 542046 471824 542096 471880
rect 542004 471822 542096 471824
rect 542004 471820 542051 471822
rect 541985 471819 542051 471820
rect 544142 471474 544148 471476
rect 542892 471414 544148 471474
rect 544142 471412 544148 471414
rect 544212 471412 544218 471476
rect 579981 470114 580047 470117
rect 583520 470114 584960 470204
rect 579981 470112 584960 470114
rect 579981 470056 579986 470112
rect 580042 470056 584960 470112
rect 579981 470054 584960 470056
rect 579981 470051 580047 470054
rect 583520 469964 584960 470054
rect 541750 468284 541756 468348
rect 541820 468284 541826 468348
rect 541758 468076 541818 468284
rect 541750 468012 541756 468076
rect 541820 468012 541826 468076
rect -960 467394 480 467484
rect 3141 467394 3207 467397
rect -960 467392 3207 467394
rect -960 467336 3146 467392
rect 3202 467336 3207 467392
rect -960 467334 3207 467336
rect -960 467244 480 467334
rect 3141 467331 3207 467334
rect 39297 467258 39363 467261
rect 39297 467256 41124 467258
rect 39297 467200 39302 467256
rect 39358 467200 41124 467256
rect 39297 467198 41124 467200
rect 39297 467195 39363 467198
rect 544653 466850 544719 466853
rect 542892 466848 544719 466850
rect 542892 466792 544658 466848
rect 544714 466792 544719 466848
rect 542892 466790 544719 466792
rect 544653 466787 544719 466790
rect 541985 466308 542051 466309
rect 541934 466306 541940 466308
rect 541894 466246 541940 466306
rect 542004 466304 542051 466308
rect 542046 466248 542051 466304
rect 541934 466244 541940 466246
rect 542004 466244 542051 466248
rect 541985 466243 542051 466244
rect 580533 465218 580599 465221
rect 583520 465218 584960 465308
rect 580533 465216 584960 465218
rect 580533 465160 580538 465216
rect 580594 465160 584960 465216
rect 580533 465158 584960 465160
rect 580533 465155 580599 465158
rect 583520 465068 584960 465158
rect 38745 462906 38811 462909
rect 38745 462904 41124 462906
rect 38745 462848 38750 462904
rect 38806 462848 41124 462904
rect 38745 462846 41124 462848
rect 38745 462843 38811 462846
rect 544653 462634 544719 462637
rect 542892 462632 544719 462634
rect -960 462498 480 462588
rect 542892 462576 544658 462632
rect 544714 462576 544719 462632
rect 542892 462574 544719 462576
rect 544653 462571 544719 462574
rect 3141 462498 3207 462501
rect -960 462496 3207 462498
rect -960 462440 3146 462496
rect 3202 462440 3207 462496
rect -960 462438 3207 462440
rect -960 462348 480 462438
rect 3141 462435 3207 462438
rect 580165 460322 580231 460325
rect 583520 460322 584960 460412
rect 580165 460320 584960 460322
rect 580165 460264 580170 460320
rect 580226 460264 584960 460320
rect 580165 460262 584960 460264
rect 580165 460259 580231 460262
rect 583520 460172 584960 460262
rect 38745 458282 38811 458285
rect 543917 458282 543983 458285
rect 38745 458280 41124 458282
rect 38745 458224 38750 458280
rect 38806 458224 41124 458280
rect 38745 458222 41124 458224
rect 542892 458280 543983 458282
rect 542892 458224 543922 458280
rect 543978 458224 543983 458280
rect 542892 458222 543983 458224
rect 38745 458219 38811 458222
rect 543917 458219 543983 458222
rect -960 457602 480 457692
rect 3233 457602 3299 457605
rect -960 457600 3299 457602
rect -960 457544 3238 457600
rect 3294 457544 3299 457600
rect -960 457542 3299 457544
rect -960 457452 480 457542
rect 3233 457539 3299 457542
rect 580165 455426 580231 455429
rect 583520 455426 584960 455516
rect 580165 455424 584960 455426
rect 580165 455368 580170 455424
rect 580226 455368 584960 455424
rect 580165 455366 584960 455368
rect 580165 455363 580231 455366
rect 583520 455276 584960 455366
rect 39481 453930 39547 453933
rect 39481 453928 41124 453930
rect 39481 453872 39486 453928
rect 39542 453872 41124 453928
rect 39481 453870 41124 453872
rect 39481 453867 39547 453870
rect 544653 453522 544719 453525
rect 542892 453520 544719 453522
rect 542892 453464 544658 453520
rect 544714 453464 544719 453520
rect 542892 453462 544719 453464
rect 544653 453459 544719 453462
rect -960 452706 480 452796
rect 3233 452706 3299 452709
rect -960 452704 3299 452706
rect -960 452648 3238 452704
rect 3294 452648 3299 452704
rect -960 452646 3299 452648
rect -960 452556 480 452646
rect 3233 452643 3299 452646
rect 580165 450530 580231 450533
rect 583520 450530 584960 450620
rect 580165 450528 584960 450530
rect 580165 450472 580170 450528
rect 580226 450472 584960 450528
rect 580165 450470 584960 450472
rect 580165 450467 580231 450470
rect 583520 450380 584960 450470
rect 39941 449306 40007 449309
rect 544653 449306 544719 449309
rect 39941 449304 41124 449306
rect 39941 449248 39946 449304
rect 40002 449248 41124 449304
rect 39941 449246 41124 449248
rect 542892 449304 544719 449306
rect 542892 449248 544658 449304
rect 544714 449248 544719 449304
rect 542892 449246 544719 449248
rect 39941 449243 40007 449246
rect 544653 449243 544719 449246
rect -960 447810 480 447900
rect 3141 447810 3207 447813
rect -960 447808 3207 447810
rect -960 447752 3146 447808
rect 3202 447752 3207 447808
rect -960 447750 3207 447752
rect -960 447660 480 447750
rect 3141 447747 3207 447750
rect 541934 445708 541940 445772
rect 542004 445770 542010 445772
rect 544653 445770 544719 445773
rect 542004 445768 544719 445770
rect 542004 445712 544658 445768
rect 544714 445712 544719 445768
rect 542004 445710 544719 445712
rect 542004 445708 542010 445710
rect 544653 445707 544719 445710
rect 580165 445634 580231 445637
rect 583520 445634 584960 445724
rect 580165 445632 584960 445634
rect 580165 445576 580170 445632
rect 580226 445576 584960 445632
rect 580165 445574 584960 445576
rect 580165 445571 580231 445574
rect 583520 445484 584960 445574
rect 38745 444818 38811 444821
rect 38745 444816 41124 444818
rect 38745 444760 38750 444816
rect 38806 444760 41124 444816
rect 38745 444758 41124 444760
rect 38745 444755 38811 444758
rect 541758 444412 541818 444516
rect 541750 444348 541756 444412
rect 541820 444348 541826 444412
rect -960 442914 480 443004
rect 3233 442914 3299 442917
rect -960 442912 3299 442914
rect -960 442856 3238 442912
rect 3294 442856 3299 442912
rect -960 442854 3299 442856
rect -960 442764 480 442854
rect 3233 442851 3299 442854
rect 541750 442444 541756 442508
rect 541820 442506 541826 442508
rect 541985 442506 542051 442509
rect 541820 442504 542051 442506
rect 541820 442448 541990 442504
rect 542046 442448 542051 442504
rect 541820 442446 542051 442448
rect 541820 442444 541826 442446
rect 541985 442443 542051 442446
rect 580165 440738 580231 440741
rect 583520 440738 584960 440828
rect 580165 440736 584960 440738
rect 580165 440680 580170 440736
rect 580226 440680 584960 440736
rect 580165 440678 584960 440680
rect 580165 440675 580231 440678
rect 583520 440588 584960 440678
rect 40217 440466 40283 440469
rect 40217 440464 41124 440466
rect 40217 440408 40222 440464
rect 40278 440408 41124 440464
rect 40217 440406 41124 440408
rect 40217 440403 40283 440406
rect 544929 440330 544995 440333
rect 542892 440328 544995 440330
rect 542892 440272 544934 440328
rect 544990 440272 544995 440328
rect 542892 440270 544995 440272
rect 544929 440267 544995 440270
rect 541750 439044 541756 439108
rect 541820 439106 541826 439108
rect 542077 439106 542143 439109
rect 541820 439104 542143 439106
rect 541820 439048 542082 439104
rect 542138 439048 542143 439104
rect 541820 439046 542143 439048
rect 541820 439044 541826 439046
rect 542077 439043 542143 439046
rect 541750 438908 541756 438972
rect 541820 438970 541826 438972
rect 541985 438970 542051 438973
rect 541820 438968 542051 438970
rect 541820 438912 541990 438968
rect 542046 438912 542051 438968
rect 541820 438910 542051 438912
rect 541820 438908 541826 438910
rect 541985 438907 542051 438910
rect -960 438018 480 438108
rect 541750 438092 541756 438156
rect 541820 438154 541826 438156
rect 542077 438154 542143 438157
rect 541820 438152 542143 438154
rect 541820 438096 542082 438152
rect 542138 438096 542143 438152
rect 541820 438094 542143 438096
rect 541820 438092 541826 438094
rect 542077 438091 542143 438094
rect 3233 438018 3299 438021
rect -960 438016 3299 438018
rect -960 437960 3238 438016
rect 3294 437960 3299 438016
rect -960 437958 3299 437960
rect -960 437868 480 437958
rect 3233 437955 3299 437958
rect 39297 435978 39363 435981
rect 39297 435976 41124 435978
rect 39297 435920 39302 435976
rect 39358 435920 41124 435976
rect 39297 435918 41124 435920
rect 39297 435915 39363 435918
rect 580165 435842 580231 435845
rect 583520 435842 584960 435932
rect 580165 435840 584960 435842
rect 580165 435784 580170 435840
rect 580226 435784 584960 435840
rect 580165 435782 584960 435784
rect 580165 435779 580231 435782
rect 543917 435706 543983 435709
rect 542892 435704 543983 435706
rect 542892 435648 543922 435704
rect 543978 435648 543983 435704
rect 583520 435692 584960 435782
rect 542892 435646 543983 435648
rect 543917 435643 543983 435646
rect -960 433122 480 433212
rect 2957 433122 3023 433125
rect -960 433120 3023 433122
rect -960 433064 2962 433120
rect 3018 433064 3023 433120
rect -960 433062 3023 433064
rect -960 432972 480 433062
rect 2957 433059 3023 433062
rect 38745 431626 38811 431629
rect 38745 431624 41124 431626
rect 38745 431568 38750 431624
rect 38806 431568 41124 431624
rect 38745 431566 41124 431568
rect 38745 431563 38811 431566
rect 543917 431354 543983 431357
rect 542892 431352 543983 431354
rect 542892 431296 543922 431352
rect 543978 431296 543983 431352
rect 542892 431294 543983 431296
rect 543917 431291 543983 431294
rect 579613 430674 579679 430677
rect 583520 430674 584960 430764
rect 579613 430672 584960 430674
rect 579613 430616 579618 430672
rect 579674 430616 584960 430672
rect 579613 430614 584960 430616
rect 579613 430611 579679 430614
rect 583520 430524 584960 430614
rect -960 427954 480 428044
rect 3233 427954 3299 427957
rect -960 427952 3299 427954
rect -960 427896 3238 427952
rect 3294 427896 3299 427952
rect -960 427894 3299 427896
rect -960 427804 480 427894
rect 3233 427891 3299 427894
rect 38745 426866 38811 426869
rect 38745 426864 41124 426866
rect 38745 426808 38750 426864
rect 38806 426808 41124 426864
rect 38745 426806 41124 426808
rect 38745 426803 38811 426806
rect 544009 426730 544075 426733
rect 542892 426728 544075 426730
rect 542892 426672 544014 426728
rect 544070 426672 544075 426728
rect 542892 426670 544075 426672
rect 544009 426667 544075 426670
rect 580165 425778 580231 425781
rect 583520 425778 584960 425868
rect 580165 425776 584960 425778
rect 580165 425720 580170 425776
rect 580226 425720 584960 425776
rect 580165 425718 584960 425720
rect 580165 425715 580231 425718
rect 583520 425628 584960 425718
rect -960 423058 480 423148
rect 3233 423058 3299 423061
rect -960 423056 3299 423058
rect -960 423000 3238 423056
rect 3294 423000 3299 423056
rect -960 422998 3299 423000
rect -960 422908 480 422998
rect 3233 422995 3299 422998
rect 39389 422650 39455 422653
rect 39389 422648 41124 422650
rect 39389 422592 39394 422648
rect 39450 422592 41124 422648
rect 39389 422590 41124 422592
rect 39389 422587 39455 422590
rect 543273 422378 543339 422381
rect 542892 422376 543339 422378
rect 542892 422320 543278 422376
rect 543334 422320 543339 422376
rect 542892 422318 543339 422320
rect 543273 422315 543339 422318
rect 580625 420882 580691 420885
rect 583520 420882 584960 420972
rect 580625 420880 584960 420882
rect 580625 420824 580630 420880
rect 580686 420824 584960 420880
rect 580625 420822 584960 420824
rect 580625 420819 580691 420822
rect 583520 420732 584960 420822
rect -960 418162 480 418252
rect 3233 418162 3299 418165
rect -960 418160 3299 418162
rect -960 418104 3238 418160
rect 3294 418104 3299 418160
rect -960 418102 3299 418104
rect -960 418012 480 418102
rect 3233 418099 3299 418102
rect 40861 418026 40927 418029
rect 40861 418024 41124 418026
rect 40861 417968 40866 418024
rect 40922 417968 41124 418024
rect 40861 417966 41124 417968
rect 40861 417963 40927 417966
rect 544193 417754 544259 417757
rect 542892 417752 544259 417754
rect 542892 417696 544198 417752
rect 544254 417696 544259 417752
rect 542892 417694 544259 417696
rect 544193 417691 544259 417694
rect 580533 415986 580599 415989
rect 583520 415986 584960 416076
rect 580533 415984 584960 415986
rect 580533 415928 580538 415984
rect 580594 415928 584960 415984
rect 580533 415926 584960 415928
rect 580533 415923 580599 415926
rect 583520 415836 584960 415926
rect 38745 413538 38811 413541
rect 38745 413536 41124 413538
rect 38745 413480 38750 413536
rect 38806 413480 41124 413536
rect 38745 413478 41124 413480
rect 38745 413475 38811 413478
rect -960 413266 480 413356
rect 3141 413266 3207 413269
rect 543917 413266 543983 413269
rect -960 413264 3207 413266
rect -960 413208 3146 413264
rect 3202 413208 3207 413264
rect -960 413206 3207 413208
rect 542892 413264 543983 413266
rect 542892 413208 543922 413264
rect 543978 413208 543983 413264
rect 542892 413206 543983 413208
rect -960 413116 480 413206
rect 3141 413203 3207 413206
rect 543917 413203 543983 413206
rect 580165 411090 580231 411093
rect 583520 411090 584960 411180
rect 580165 411088 584960 411090
rect 580165 411032 580170 411088
rect 580226 411032 584960 411088
rect 580165 411030 584960 411032
rect 580165 411027 580231 411030
rect 583520 410940 584960 411030
rect 40769 409050 40835 409053
rect 40769 409048 41124 409050
rect 40769 408992 40774 409048
rect 40830 408992 41124 409048
rect 40769 408990 41124 408992
rect 40769 408987 40835 408990
rect 544193 408778 544259 408781
rect 542892 408776 544259 408778
rect 542892 408720 544198 408776
rect 544254 408720 544259 408776
rect 542892 408718 544259 408720
rect 544193 408715 544259 408718
rect -960 408370 480 408460
rect 2773 408370 2839 408373
rect -960 408368 2839 408370
rect -960 408312 2778 408368
rect 2834 408312 2839 408368
rect -960 408310 2839 408312
rect -960 408220 480 408310
rect 2773 408307 2839 408310
rect 580165 406194 580231 406197
rect 583520 406194 584960 406284
rect 580165 406192 584960 406194
rect 580165 406136 580170 406192
rect 580226 406136 584960 406192
rect 580165 406134 584960 406136
rect 580165 406131 580231 406134
rect 583520 406044 584960 406134
rect 40166 404500 40172 404564
rect 40236 404562 40242 404564
rect 40236 404502 41124 404562
rect 40236 404500 40242 404502
rect 544929 404426 544995 404429
rect 542892 404424 544995 404426
rect 542892 404368 544934 404424
rect 544990 404368 544995 404424
rect 542892 404366 544995 404368
rect 544929 404363 544995 404366
rect -960 403474 480 403564
rect 3233 403474 3299 403477
rect -960 403472 3299 403474
rect -960 403416 3238 403472
rect 3294 403416 3299 403472
rect -960 403414 3299 403416
rect -960 403324 480 403414
rect 3233 403411 3299 403414
rect 579705 401298 579771 401301
rect 583520 401298 584960 401388
rect 579705 401296 584960 401298
rect 579705 401240 579710 401296
rect 579766 401240 584960 401296
rect 579705 401238 584960 401240
rect 579705 401235 579771 401238
rect 583520 401148 584960 401238
rect 544745 400074 544811 400077
rect 542892 400072 544811 400074
rect 542892 400016 544750 400072
rect 544806 400016 544811 400072
rect 542892 400014 544811 400016
rect 544745 400011 544811 400014
rect 38745 399938 38811 399941
rect 38745 399936 41124 399938
rect 38745 399880 38750 399936
rect 38806 399880 41124 399936
rect 38745 399878 41124 399880
rect 38745 399875 38811 399878
rect -960 398578 480 398668
rect 3233 398578 3299 398581
rect -960 398576 3299 398578
rect -960 398520 3238 398576
rect 3294 398520 3299 398576
rect -960 398518 3299 398520
rect -960 398428 480 398518
rect 3233 398515 3299 398518
rect 580625 396402 580691 396405
rect 583520 396402 584960 396492
rect 580625 396400 584960 396402
rect 580625 396344 580630 396400
rect 580686 396344 584960 396400
rect 580625 396342 584960 396344
rect 580625 396339 580691 396342
rect 583520 396252 584960 396342
rect 39665 395722 39731 395725
rect 39665 395720 41124 395722
rect 39665 395664 39670 395720
rect 39726 395664 41124 395720
rect 39665 395662 41124 395664
rect 39665 395659 39731 395662
rect 544745 395450 544811 395453
rect 542892 395448 544811 395450
rect 542892 395392 544750 395448
rect 544806 395392 544811 395448
rect 542892 395390 544811 395392
rect 544745 395387 544811 395390
rect -960 393682 480 393772
rect 2773 393682 2839 393685
rect -960 393680 2839 393682
rect -960 393624 2778 393680
rect 2834 393624 2839 393680
rect -960 393622 2839 393624
rect -960 393532 480 393622
rect 2773 393619 2839 393622
rect 579613 391506 579679 391509
rect 583520 391506 584960 391596
rect 579613 391504 584960 391506
rect 579613 391448 579618 391504
rect 579674 391448 584960 391504
rect 579613 391446 584960 391448
rect 579613 391443 579679 391446
rect 583520 391356 584960 391446
rect 39573 391098 39639 391101
rect 39573 391096 41124 391098
rect 39573 391040 39578 391096
rect 39634 391040 41124 391096
rect 39573 391038 41124 391040
rect 39573 391035 39639 391038
rect 544745 390962 544811 390965
rect 542892 390960 544811 390962
rect 542892 390904 544750 390960
rect 544806 390904 544811 390960
rect 542892 390902 544811 390904
rect 544745 390899 544811 390902
rect -960 388786 480 388876
rect 3969 388786 4035 388789
rect -960 388784 4035 388786
rect -960 388728 3974 388784
rect 4030 388728 4035 388784
rect -960 388726 4035 388728
rect -960 388636 480 388726
rect 3969 388723 4035 388726
rect 41045 387290 41111 387293
rect 41045 387288 41154 387290
rect 41045 387232 41050 387288
rect 41106 387232 41154 387288
rect 41045 387227 41154 387232
rect 41094 386716 41154 387227
rect 580165 386610 580231 386613
rect 583520 386610 584960 386700
rect 580165 386608 584960 386610
rect 580165 386552 580170 386608
rect 580226 386552 584960 386608
rect 580165 386550 584960 386552
rect 580165 386547 580231 386550
rect 544929 386474 544995 386477
rect 542892 386472 544995 386474
rect 542892 386416 544934 386472
rect 544990 386416 544995 386472
rect 583520 386460 584960 386550
rect 542892 386414 544995 386416
rect 544929 386411 544995 386414
rect -960 383890 480 383980
rect 2773 383890 2839 383893
rect -960 383888 2839 383890
rect -960 383832 2778 383888
rect 2834 383832 2839 383888
rect -960 383830 2839 383832
rect -960 383740 480 383830
rect 2773 383827 2839 383830
rect 39062 382332 39068 382396
rect 39132 382394 39138 382396
rect 39132 382334 41124 382394
rect 39132 382332 39138 382334
rect 544193 381986 544259 381989
rect 542892 381984 544259 381986
rect 542892 381928 544198 381984
rect 544254 381928 544259 381984
rect 542892 381926 544259 381928
rect 544193 381923 544259 381926
rect 579797 381714 579863 381717
rect 583520 381714 584960 381804
rect 579797 381712 584960 381714
rect 579797 381656 579802 381712
rect 579858 381656 584960 381712
rect 579797 381654 584960 381656
rect 579797 381651 579863 381654
rect 583520 381564 584960 381654
rect -960 378844 480 379084
rect 39389 377770 39455 377773
rect 39389 377768 41124 377770
rect 39389 377712 39394 377768
rect 39450 377712 41124 377768
rect 39389 377710 41124 377712
rect 39389 377707 39455 377710
rect 544745 377498 544811 377501
rect 542892 377496 544811 377498
rect 542892 377440 544750 377496
rect 544806 377440 544811 377496
rect 542892 377438 544811 377440
rect 544745 377435 544811 377438
rect 580165 376546 580231 376549
rect 583520 376546 584960 376636
rect 580165 376544 584960 376546
rect 580165 376488 580170 376544
rect 580226 376488 584960 376544
rect 580165 376486 584960 376488
rect 580165 376483 580231 376486
rect 583520 376396 584960 376486
rect -960 373826 480 373916
rect 3969 373826 4035 373829
rect -960 373824 4035 373826
rect -960 373768 3974 373824
rect 4030 373768 4035 373824
rect -960 373766 4035 373768
rect -960 373676 480 373766
rect 3969 373763 4035 373766
rect 39389 373282 39455 373285
rect 39389 373280 41124 373282
rect 39389 373224 39394 373280
rect 39450 373224 41124 373280
rect 39389 373222 41124 373224
rect 39389 373219 39455 373222
rect 544009 373010 544075 373013
rect 542892 373008 544075 373010
rect 542892 372952 544014 373008
rect 544070 372952 544075 373008
rect 542892 372950 544075 372952
rect 544009 372947 544075 372950
rect 579613 371650 579679 371653
rect 583520 371650 584960 371740
rect 579613 371648 584960 371650
rect 579613 371592 579618 371648
rect 579674 371592 584960 371648
rect 579613 371590 584960 371592
rect 579613 371587 579679 371590
rect 583520 371500 584960 371590
rect 543038 369140 543044 369204
rect 543108 369202 543114 369204
rect 544101 369202 544167 369205
rect 543108 369200 544167 369202
rect 543108 369144 544106 369200
rect 544162 369144 544167 369200
rect 543108 369142 544167 369144
rect 543108 369140 543114 369142
rect 544101 369139 544167 369142
rect -960 368930 480 369020
rect 3233 368930 3299 368933
rect -960 368928 3299 368930
rect -960 368872 3238 368928
rect 3294 368872 3299 368928
rect -960 368870 3299 368872
rect -960 368780 480 368870
rect 3233 368867 3299 368870
rect 39573 368658 39639 368661
rect 39573 368656 41124 368658
rect 39573 368600 39578 368656
rect 39634 368600 41124 368656
rect 39573 368598 41124 368600
rect 39573 368595 39639 368598
rect 544101 368522 544167 368525
rect 542892 368520 544167 368522
rect 542892 368464 544106 368520
rect 544162 368464 544167 368520
rect 542892 368462 544167 368464
rect 544101 368459 544167 368462
rect 580165 366754 580231 366757
rect 583520 366754 584960 366844
rect 580165 366752 584960 366754
rect 580165 366696 580170 366752
rect 580226 366696 584960 366752
rect 580165 366694 584960 366696
rect 580165 366691 580231 366694
rect 583520 366604 584960 366694
rect 39062 364380 39068 364444
rect 39132 364442 39138 364444
rect 39132 364382 41124 364442
rect 39132 364380 39138 364382
rect 544745 364170 544811 364173
rect 542892 364168 544811 364170
rect -960 364034 480 364124
rect 542892 364112 544750 364168
rect 544806 364112 544811 364168
rect 542892 364110 544811 364112
rect 544745 364107 544811 364110
rect 3325 364034 3391 364037
rect -960 364032 3391 364034
rect -960 363976 3330 364032
rect 3386 363976 3391 364032
rect -960 363974 3391 363976
rect -960 363884 480 363974
rect 3325 363971 3391 363974
rect 580165 361858 580231 361861
rect 583520 361858 584960 361948
rect 580165 361856 584960 361858
rect 580165 361800 580170 361856
rect 580226 361800 584960 361856
rect 580165 361798 584960 361800
rect 580165 361795 580231 361798
rect 583520 361708 584960 361798
rect 38878 359756 38884 359820
rect 38948 359818 38954 359820
rect 38948 359758 41124 359818
rect 38948 359756 38954 359758
rect 544929 359410 544995 359413
rect 542892 359408 544995 359410
rect 542892 359352 544934 359408
rect 544990 359352 544995 359408
rect 542892 359350 544995 359352
rect 544929 359347 544995 359350
rect -960 359138 480 359228
rect 4061 359138 4127 359141
rect -960 359136 4127 359138
rect -960 359080 4066 359136
rect 4122 359080 4127 359136
rect -960 359078 4127 359080
rect -960 358988 480 359078
rect 4061 359075 4127 359078
rect 579981 356962 580047 356965
rect 583520 356962 584960 357052
rect 579981 356960 584960 356962
rect 579981 356904 579986 356960
rect 580042 356904 584960 356960
rect 579981 356902 584960 356904
rect 579981 356899 580047 356902
rect 583520 356812 584960 356902
rect 40953 356010 41019 356013
rect 40953 356008 41154 356010
rect 40953 355952 40958 356008
rect 41014 355952 41154 356008
rect 40953 355950 41154 355952
rect 40953 355947 41019 355950
rect 41094 355436 41154 355950
rect 543089 355194 543155 355197
rect 542892 355192 543155 355194
rect 542892 355136 543094 355192
rect 543150 355136 543155 355192
rect 542892 355134 543155 355136
rect 543089 355131 543155 355134
rect -960 354242 480 354332
rect 3141 354242 3207 354245
rect -960 354240 3207 354242
rect -960 354184 3146 354240
rect 3202 354184 3207 354240
rect -960 354182 3207 354184
rect -960 354092 480 354182
rect 3141 354179 3207 354182
rect 580165 352066 580231 352069
rect 583520 352066 584960 352156
rect 580165 352064 584960 352066
rect 580165 352008 580170 352064
rect 580226 352008 584960 352064
rect 580165 352006 584960 352008
rect 580165 352003 580231 352006
rect 583520 351916 584960 352006
rect 38745 350706 38811 350709
rect 38745 350704 41124 350706
rect 38745 350648 38750 350704
rect 38806 350648 41124 350704
rect 38745 350646 41124 350648
rect 38745 350643 38811 350646
rect 542862 350301 542922 350404
rect 542862 350296 542971 350301
rect 542862 350240 542910 350296
rect 542966 350240 542971 350296
rect 542862 350238 542971 350240
rect 542905 350235 542971 350238
rect -960 349346 480 349436
rect 2773 349346 2839 349349
rect -960 349344 2839 349346
rect -960 349288 2778 349344
rect 2834 349288 2839 349344
rect -960 349286 2839 349288
rect -960 349196 480 349286
rect 2773 349283 2839 349286
rect 580165 347170 580231 347173
rect 583520 347170 584960 347260
rect 580165 347168 584960 347170
rect 580165 347112 580170 347168
rect 580226 347112 584960 347168
rect 580165 347110 584960 347112
rect 580165 347107 580231 347110
rect 583520 347020 584960 347110
rect 38745 346490 38811 346493
rect 38745 346488 41124 346490
rect 38745 346432 38750 346488
rect 38806 346432 41124 346488
rect 38745 346430 41124 346432
rect 38745 346427 38811 346430
rect 544561 346218 544627 346221
rect 542892 346216 544627 346218
rect 542892 346160 544566 346216
rect 544622 346160 544627 346216
rect 542892 346158 544627 346160
rect 544561 346155 544627 346158
rect -960 344450 480 344540
rect 3325 344450 3391 344453
rect -960 344448 3391 344450
rect -960 344392 3330 344448
rect 3386 344392 3391 344448
rect -960 344390 3391 344392
rect -960 344300 480 344390
rect 3325 344387 3391 344390
rect 580717 342274 580783 342277
rect 583520 342274 584960 342364
rect 580717 342272 584960 342274
rect 580717 342216 580722 342272
rect 580778 342216 584960 342272
rect 580717 342214 584960 342216
rect 580717 342211 580783 342214
rect 583520 342124 584960 342214
rect 544745 341866 544811 341869
rect 542892 341864 544811 341866
rect 542892 341808 544750 341864
rect 544806 341808 544811 341864
rect 542892 341806 544811 341808
rect 544745 341803 544811 341806
rect 39665 341730 39731 341733
rect 39665 341728 41124 341730
rect 39665 341672 39670 341728
rect 39726 341672 41124 341728
rect 39665 341670 41124 341672
rect 39665 341667 39731 341670
rect -960 339554 480 339644
rect 3325 339554 3391 339557
rect -960 339552 3391 339554
rect -960 339496 3330 339552
rect 3386 339496 3391 339552
rect -960 339494 3391 339496
rect -960 339404 480 339494
rect 3325 339491 3391 339494
rect 38878 337316 38884 337380
rect 38948 337378 38954 337380
rect 580165 337378 580231 337381
rect 583520 337378 584960 337468
rect 38948 337318 41124 337378
rect 580165 337376 584960 337378
rect 580165 337320 580170 337376
rect 580226 337320 584960 337376
rect 580165 337318 584960 337320
rect 38948 337316 38954 337318
rect 580165 337315 580231 337318
rect 583520 337228 584960 337318
rect 544561 337106 544627 337109
rect 542892 337104 544627 337106
rect 542892 337048 544566 337104
rect 544622 337048 544627 337104
rect 542892 337046 544627 337048
rect 544561 337043 544627 337046
rect -960 334658 480 334748
rect 2957 334658 3023 334661
rect -960 334656 3023 334658
rect -960 334600 2962 334656
rect 3018 334600 3023 334656
rect -960 334598 3023 334600
rect -960 334508 480 334598
rect 2957 334595 3023 334598
rect 544469 332890 544535 332893
rect 542892 332888 544535 332890
rect 542892 332832 544474 332888
rect 544530 332832 544535 332888
rect 542892 332830 544535 332832
rect 544469 332827 544535 332830
rect 38745 332754 38811 332757
rect 38745 332752 41124 332754
rect 38745 332696 38750 332752
rect 38806 332696 41124 332752
rect 38745 332694 41124 332696
rect 38745 332691 38811 332694
rect 580717 332482 580783 332485
rect 583520 332482 584960 332572
rect 580717 332480 584960 332482
rect 580717 332424 580722 332480
rect 580778 332424 584960 332480
rect 580717 332422 584960 332424
rect 580717 332419 580783 332422
rect 583520 332332 584960 332422
rect -960 329762 480 329852
rect 3233 329762 3299 329765
rect -960 329760 3299 329762
rect -960 329704 3238 329760
rect 3294 329704 3299 329760
rect -960 329702 3299 329704
rect -960 329612 480 329702
rect 3233 329699 3299 329702
rect 40585 328538 40651 328541
rect 40585 328536 41124 328538
rect 40585 328480 40590 328536
rect 40646 328480 41124 328536
rect 40585 328478 41124 328480
rect 40585 328475 40651 328478
rect 544377 328266 544443 328269
rect 542892 328264 544443 328266
rect 542892 328208 544382 328264
rect 544438 328208 544443 328264
rect 542892 328206 544443 328208
rect 544377 328203 544443 328206
rect 579981 327586 580047 327589
rect 583520 327586 584960 327676
rect 579981 327584 584960 327586
rect 579981 327528 579986 327584
rect 580042 327528 584960 327584
rect 579981 327526 584960 327528
rect 579981 327523 580047 327526
rect 583520 327436 584960 327526
rect -960 324866 480 324956
rect 4061 324866 4127 324869
rect -960 324864 4127 324866
rect -960 324808 4066 324864
rect 4122 324808 4127 324864
rect -960 324806 4127 324808
rect -960 324716 480 324806
rect 4061 324803 4127 324806
rect 38745 324186 38811 324189
rect 38745 324184 41124 324186
rect 38745 324128 38750 324184
rect 38806 324128 41124 324184
rect 38745 324126 41124 324128
rect 38745 324123 38811 324126
rect 544285 323914 544351 323917
rect 542892 323912 544351 323914
rect 542892 323856 544290 323912
rect 544346 323856 544351 323912
rect 542892 323854 544351 323856
rect 544285 323851 544351 323854
rect 579797 322418 579863 322421
rect 583520 322418 584960 322508
rect 579797 322416 584960 322418
rect 579797 322360 579802 322416
rect 579858 322360 584960 322416
rect 579797 322358 584960 322360
rect 579797 322355 579863 322358
rect 583520 322268 584960 322358
rect -960 319698 480 319788
rect 3325 319698 3391 319701
rect -960 319696 3391 319698
rect -960 319640 3330 319696
rect 3386 319640 3391 319696
rect -960 319638 3391 319640
rect -960 319548 480 319638
rect 3325 319635 3391 319638
rect 39297 319426 39363 319429
rect 39297 319424 41124 319426
rect 39297 319368 39302 319424
rect 39358 319368 41124 319424
rect 39297 319366 41124 319368
rect 39297 319363 39363 319366
rect 544929 319154 544995 319157
rect 542892 319152 544995 319154
rect 542892 319096 544934 319152
rect 544990 319096 544995 319152
rect 542892 319094 544995 319096
rect 544929 319091 544995 319094
rect 580809 317522 580875 317525
rect 583520 317522 584960 317612
rect 580809 317520 584960 317522
rect 580809 317464 580814 317520
rect 580870 317464 584960 317520
rect 580809 317462 584960 317464
rect 580809 317459 580875 317462
rect 583520 317372 584960 317462
rect 38745 315074 38811 315077
rect 38745 315072 41124 315074
rect 38745 315016 38750 315072
rect 38806 315016 41124 315072
rect 38745 315014 41124 315016
rect 38745 315011 38811 315014
rect -960 314802 480 314892
rect 3325 314802 3391 314805
rect 544285 314802 544351 314805
rect -960 314800 3391 314802
rect -960 314744 3330 314800
rect 3386 314744 3391 314800
rect -960 314742 3391 314744
rect 542892 314800 544351 314802
rect 542892 314744 544290 314800
rect 544346 314744 544351 314800
rect 542892 314742 544351 314744
rect -960 314652 480 314742
rect 3325 314739 3391 314742
rect 544285 314739 544351 314742
rect 580165 312626 580231 312629
rect 583520 312626 584960 312716
rect 580165 312624 584960 312626
rect 580165 312568 580170 312624
rect 580226 312568 584960 312624
rect 580165 312566 584960 312568
rect 580165 312563 580231 312566
rect 583520 312476 584960 312566
rect 38745 310586 38811 310589
rect 38745 310584 41124 310586
rect 38745 310528 38750 310584
rect 38806 310528 41124 310584
rect 38745 310526 41124 310528
rect 38745 310523 38811 310526
rect 544377 310178 544443 310181
rect 542892 310176 544443 310178
rect 542892 310120 544382 310176
rect 544438 310120 544443 310176
rect 542892 310118 544443 310120
rect 544377 310115 544443 310118
rect -960 309906 480 309996
rect 2957 309906 3023 309909
rect -960 309904 3023 309906
rect -960 309848 2962 309904
rect 3018 309848 3023 309904
rect -960 309846 3023 309848
rect -960 309756 480 309846
rect 2957 309843 3023 309846
rect 580165 307730 580231 307733
rect 583520 307730 584960 307820
rect 580165 307728 584960 307730
rect 580165 307672 580170 307728
rect 580226 307672 584960 307728
rect 580165 307670 584960 307672
rect 580165 307667 580231 307670
rect 583520 307580 584960 307670
rect 38745 306234 38811 306237
rect 38745 306232 41124 306234
rect 38745 306176 38750 306232
rect 38806 306176 41124 306232
rect 38745 306174 41124 306176
rect 38745 306171 38811 306174
rect 542862 305285 542922 305796
rect 542862 305280 542971 305285
rect 542862 305224 542910 305280
rect 542966 305224 542971 305280
rect 542862 305222 542971 305224
rect 542905 305219 542971 305222
rect -960 305010 480 305100
rect 2773 305010 2839 305013
rect -960 305008 2839 305010
rect -960 304952 2778 305008
rect 2834 304952 2839 305008
rect -960 304950 2839 304952
rect -960 304860 480 304950
rect 2773 304947 2839 304950
rect 580165 302834 580231 302837
rect 583520 302834 584960 302924
rect 580165 302832 584960 302834
rect 580165 302776 580170 302832
rect 580226 302776 584960 302832
rect 580165 302774 584960 302776
rect 580165 302771 580231 302774
rect 583520 302684 584960 302774
rect 542813 301882 542879 301885
rect 542813 301880 542922 301882
rect 542813 301824 542818 301880
rect 542874 301824 542922 301880
rect 542813 301819 542922 301824
rect 40401 301610 40467 301613
rect 40401 301608 41124 301610
rect 40401 301552 40406 301608
rect 40462 301552 41124 301608
rect 40401 301550 41124 301552
rect 40401 301547 40467 301550
rect 542862 301308 542922 301819
rect -960 300114 480 300204
rect 3325 300114 3391 300117
rect -960 300112 3391 300114
rect -960 300056 3330 300112
rect 3386 300056 3391 300112
rect -960 300054 3391 300056
rect -960 299964 480 300054
rect 3325 300051 3391 300054
rect 579613 297938 579679 297941
rect 583520 297938 584960 298028
rect 579613 297936 584960 297938
rect 579613 297880 579618 297936
rect 579674 297880 584960 297936
rect 579613 297878 584960 297880
rect 579613 297875 579679 297878
rect 583520 297788 584960 297878
rect 40401 297122 40467 297125
rect 40401 297120 41124 297122
rect 40401 297064 40406 297120
rect 40462 297064 41124 297120
rect 40401 297062 41124 297064
rect 40401 297059 40467 297062
rect 542678 296716 542738 296820
rect 542670 296652 542676 296716
rect 542740 296652 542746 296716
rect -960 295218 480 295308
rect 3325 295218 3391 295221
rect -960 295216 3391 295218
rect -960 295160 3330 295216
rect 3386 295160 3391 295216
rect -960 295158 3391 295160
rect -960 295068 480 295158
rect 3325 295155 3391 295158
rect 579797 293042 579863 293045
rect 583520 293042 584960 293132
rect 579797 293040 584960 293042
rect 579797 292984 579802 293040
rect 579858 292984 584960 293040
rect 579797 292982 584960 292984
rect 579797 292979 579863 292982
rect 583520 292892 584960 292982
rect 38745 292634 38811 292637
rect 38745 292632 41124 292634
rect 38745 292576 38750 292632
rect 38806 292576 41124 292632
rect 38745 292574 41124 292576
rect 38745 292571 38811 292574
rect 542862 291685 542922 292196
rect 542813 291680 542922 291685
rect 542813 291624 542818 291680
rect 542874 291624 542922 291680
rect 542813 291622 542922 291624
rect 542813 291619 542879 291622
rect 541750 291076 541756 291140
rect 541820 291138 541826 291140
rect 547045 291138 547111 291141
rect 541820 291136 547111 291138
rect 541820 291080 547050 291136
rect 547106 291080 547111 291136
rect 541820 291078 547111 291080
rect 541820 291076 541826 291078
rect 547045 291075 547111 291078
rect -960 290322 480 290412
rect 3141 290322 3207 290325
rect -960 290320 3207 290322
rect -960 290264 3146 290320
rect 3202 290264 3207 290320
rect -960 290262 3207 290264
rect -960 290172 480 290262
rect 3141 290259 3207 290262
rect 39573 288146 39639 288149
rect 579613 288146 579679 288149
rect 583520 288146 584960 288236
rect 39573 288144 41124 288146
rect 39573 288088 39578 288144
rect 39634 288088 41124 288144
rect 39573 288086 41124 288088
rect 579613 288144 584960 288146
rect 579613 288088 579618 288144
rect 579674 288088 584960 288144
rect 579613 288086 584960 288088
rect 39573 288083 39639 288086
rect 579613 288083 579679 288086
rect 583520 287996 584960 288086
rect 545665 287874 545731 287877
rect 542892 287872 545731 287874
rect 542892 287816 545670 287872
rect 545726 287816 545731 287872
rect 542892 287814 545731 287816
rect 545665 287811 545731 287814
rect -960 285426 480 285516
rect 3233 285426 3299 285429
rect -960 285424 3299 285426
rect -960 285368 3238 285424
rect 3294 285368 3299 285424
rect -960 285366 3299 285368
rect -960 285276 480 285366
rect 3233 285363 3299 285366
rect 542486 284140 542492 284204
rect 542556 284140 542562 284204
rect 38745 283658 38811 283661
rect 38745 283656 41124 283658
rect 38745 283600 38750 283656
rect 38806 283600 41124 283656
rect 542494 283628 542554 284140
rect 38745 283598 41124 283600
rect 38745 283595 38811 283598
rect 579613 283250 579679 283253
rect 583520 283250 584960 283340
rect 579613 283248 584960 283250
rect 579613 283192 579618 283248
rect 579674 283192 584960 283248
rect 579613 283190 584960 283192
rect 579613 283187 579679 283190
rect 583520 283100 584960 283190
rect -960 280530 480 280620
rect 3325 280530 3391 280533
rect -960 280528 3391 280530
rect -960 280472 3330 280528
rect 3386 280472 3391 280528
rect -960 280470 3391 280472
rect -960 280380 480 280470
rect 3325 280467 3391 280470
rect 39297 279306 39363 279309
rect 39297 279304 41124 279306
rect 39297 279248 39302 279304
rect 39358 279248 41124 279304
rect 39297 279246 41124 279248
rect 39297 279243 39363 279246
rect 544929 278898 544995 278901
rect 542892 278896 544995 278898
rect 542892 278840 544934 278896
rect 544990 278840 544995 278896
rect 542892 278838 544995 278840
rect 544929 278835 544995 278838
rect 579981 278354 580047 278357
rect 583520 278354 584960 278444
rect 579981 278352 584960 278354
rect 579981 278296 579986 278352
rect 580042 278296 584960 278352
rect 579981 278294 584960 278296
rect 579981 278291 580047 278294
rect 583520 278204 584960 278294
rect -960 275634 480 275724
rect 3325 275634 3391 275637
rect -960 275632 3391 275634
rect -960 275576 3330 275632
rect 3386 275576 3391 275632
rect -960 275574 3391 275576
rect -960 275484 480 275574
rect 3325 275571 3391 275574
rect 40493 274682 40559 274685
rect 544745 274682 544811 274685
rect 40493 274680 41124 274682
rect 40493 274624 40498 274680
rect 40554 274624 41124 274680
rect 40493 274622 41124 274624
rect 542892 274680 544811 274682
rect 542892 274624 544750 274680
rect 544806 274624 544811 274680
rect 542892 274622 544811 274624
rect 40493 274619 40559 274622
rect 544745 274619 544811 274622
rect 580165 273458 580231 273461
rect 583520 273458 584960 273548
rect 580165 273456 584960 273458
rect 580165 273400 580170 273456
rect 580226 273400 584960 273456
rect 580165 273398 584960 273400
rect 580165 273395 580231 273398
rect 583520 273308 584960 273398
rect -960 270738 480 270828
rect 3325 270738 3391 270741
rect -960 270736 3391 270738
rect -960 270680 3330 270736
rect 3386 270680 3391 270736
rect -960 270678 3391 270680
rect -960 270588 480 270678
rect 3325 270675 3391 270678
rect 38745 270330 38811 270333
rect 38745 270328 41124 270330
rect 38745 270272 38750 270328
rect 38806 270272 41124 270328
rect 38745 270270 41124 270272
rect 38745 270267 38811 270270
rect 544929 269922 544995 269925
rect 542892 269920 544995 269922
rect 542892 269864 544934 269920
rect 544990 269864 544995 269920
rect 542892 269862 544995 269864
rect 544929 269859 544995 269862
rect 580441 268290 580507 268293
rect 583520 268290 584960 268380
rect 580441 268288 584960 268290
rect 580441 268232 580446 268288
rect 580502 268232 584960 268288
rect 580441 268230 584960 268232
rect 580441 268227 580507 268230
rect 583520 268140 584960 268230
rect 39757 265978 39823 265981
rect 39757 265976 41124 265978
rect 39757 265920 39762 265976
rect 39818 265920 41124 265976
rect 39757 265918 41124 265920
rect 39757 265915 39823 265918
rect -960 265570 480 265660
rect 3141 265570 3207 265573
rect 545481 265570 545547 265573
rect -960 265568 3207 265570
rect -960 265512 3146 265568
rect 3202 265512 3207 265568
rect -960 265510 3207 265512
rect 542892 265568 545547 265570
rect 542892 265512 545486 265568
rect 545542 265512 545547 265568
rect 542892 265510 545547 265512
rect -960 265420 480 265510
rect 3141 265507 3207 265510
rect 545481 265507 545547 265510
rect 580441 263394 580507 263397
rect 583520 263394 584960 263484
rect 580441 263392 584960 263394
rect 580441 263336 580446 263392
rect 580502 263336 584960 263392
rect 580441 263334 584960 263336
rect 580441 263331 580507 263334
rect 583520 263244 584960 263334
rect 39849 261354 39915 261357
rect 39849 261352 41124 261354
rect 39849 261296 39854 261352
rect 39910 261296 41124 261352
rect 39849 261294 41124 261296
rect 39849 261291 39915 261294
rect 544510 261082 544516 261084
rect 542892 261022 544516 261082
rect 544510 261020 544516 261022
rect 544580 261020 544586 261084
rect -960 260674 480 260764
rect 3141 260674 3207 260677
rect -960 260672 3207 260674
rect -960 260616 3146 260672
rect 3202 260616 3207 260672
rect -960 260614 3207 260616
rect -960 260524 480 260614
rect 3141 260611 3207 260614
rect 580165 258498 580231 258501
rect 583520 258498 584960 258588
rect 580165 258496 584960 258498
rect 580165 258440 580170 258496
rect 580226 258440 584960 258496
rect 580165 258438 584960 258440
rect 580165 258435 580231 258438
rect 583520 258348 584960 258438
rect 40493 256866 40559 256869
rect 40493 256864 41124 256866
rect 40493 256808 40498 256864
rect 40554 256808 41124 256864
rect 40493 256806 41124 256808
rect 40493 256803 40559 256806
rect 544745 256594 544811 256597
rect 542892 256592 544811 256594
rect 542892 256536 544750 256592
rect 544806 256536 544811 256592
rect 542892 256534 544811 256536
rect 544745 256531 544811 256534
rect -960 255778 480 255868
rect 3601 255778 3667 255781
rect -960 255776 3667 255778
rect -960 255720 3606 255776
rect 3662 255720 3667 255776
rect -960 255718 3667 255720
rect -960 255628 480 255718
rect 3601 255715 3667 255718
rect 579797 253602 579863 253605
rect 583520 253602 584960 253692
rect 579797 253600 584960 253602
rect 579797 253544 579802 253600
rect 579858 253544 584960 253600
rect 579797 253542 584960 253544
rect 579797 253539 579863 253542
rect 583520 253452 584960 253542
rect 38745 252242 38811 252245
rect 38745 252240 41124 252242
rect 38745 252184 38750 252240
rect 38806 252184 41124 252240
rect 38745 252182 41124 252184
rect 38745 252179 38811 252182
rect 543825 252106 543891 252109
rect 542892 252104 543891 252106
rect 542892 252048 543830 252104
rect 543886 252048 543891 252104
rect 542892 252046 543891 252048
rect 543825 252043 543891 252046
rect -960 250882 480 250972
rect 3785 250882 3851 250885
rect -960 250880 3851 250882
rect -960 250824 3790 250880
rect 3846 250824 3851 250880
rect -960 250822 3851 250824
rect -960 250732 480 250822
rect 3785 250819 3851 250822
rect 579613 248706 579679 248709
rect 583520 248706 584960 248796
rect 579613 248704 584960 248706
rect 579613 248648 579618 248704
rect 579674 248648 584960 248704
rect 579613 248646 584960 248648
rect 579613 248643 579679 248646
rect 583520 248556 584960 248646
rect 38837 248026 38903 248029
rect 38837 248024 41124 248026
rect 38837 247968 38842 248024
rect 38898 247968 41124 248024
rect 38837 247966 41124 247968
rect 38837 247963 38903 247966
rect 544745 247618 544811 247621
rect 542892 247616 544811 247618
rect 542892 247560 544750 247616
rect 544806 247560 544811 247616
rect 542892 247558 544811 247560
rect 544745 247555 544811 247558
rect -960 245986 480 246076
rect 3601 245986 3667 245989
rect -960 245984 3667 245986
rect -960 245928 3606 245984
rect 3662 245928 3667 245984
rect -960 245926 3667 245928
rect -960 245836 480 245926
rect 3601 245923 3667 245926
rect 580349 243810 580415 243813
rect 583520 243810 584960 243900
rect 580349 243808 584960 243810
rect 580349 243752 580354 243808
rect 580410 243752 584960 243808
rect 580349 243750 584960 243752
rect 580349 243747 580415 243750
rect 583520 243660 584960 243750
rect 38745 243402 38811 243405
rect 38745 243400 41124 243402
rect 38745 243344 38750 243400
rect 38806 243344 41124 243400
rect 38745 243342 41124 243344
rect 38745 243339 38811 243342
rect 544745 242994 544811 242997
rect 542892 242992 544811 242994
rect 542892 242936 544750 242992
rect 544806 242936 544811 242992
rect 542892 242934 544811 242936
rect 544745 242931 544811 242934
rect -960 241090 480 241180
rect 3601 241090 3667 241093
rect -960 241088 3667 241090
rect -960 241032 3606 241088
rect 3662 241032 3667 241088
rect -960 241030 3667 241032
rect -960 240940 480 241030
rect 3601 241027 3667 241030
rect 38745 239050 38811 239053
rect 38745 239048 41124 239050
rect 38745 238992 38750 239048
rect 38806 238992 41124 239048
rect 38745 238990 41124 238992
rect 38745 238987 38811 238990
rect 580165 238914 580231 238917
rect 583520 238914 584960 239004
rect 580165 238912 584960 238914
rect 580165 238856 580170 238912
rect 580226 238856 584960 238912
rect 580165 238854 584960 238856
rect 580165 238851 580231 238854
rect 583520 238764 584960 238854
rect 544745 238642 544811 238645
rect 542892 238640 544811 238642
rect 542892 238584 544750 238640
rect 544806 238584 544811 238640
rect 542892 238582 544811 238584
rect 544745 238579 544811 238582
rect -960 236194 480 236284
rect 3601 236194 3667 236197
rect -960 236192 3667 236194
rect -960 236136 3606 236192
rect 3662 236136 3667 236192
rect -960 236134 3667 236136
rect -960 236044 480 236134
rect 3601 236131 3667 236134
rect 38745 234426 38811 234429
rect 38745 234424 41124 234426
rect 38745 234368 38750 234424
rect 38806 234368 41124 234424
rect 38745 234366 41124 234368
rect 38745 234363 38811 234366
rect 544326 234154 544332 234156
rect 542892 234094 544332 234154
rect 544326 234092 544332 234094
rect 544396 234092 544402 234156
rect 579981 234018 580047 234021
rect 583520 234018 584960 234108
rect 579981 234016 584960 234018
rect 579981 233960 579986 234016
rect 580042 233960 584960 234016
rect 579981 233958 584960 233960
rect 579981 233955 580047 233958
rect 583520 233868 584960 233958
rect -960 231298 480 231388
rect 3877 231298 3943 231301
rect -960 231296 3943 231298
rect -960 231240 3882 231296
rect 3938 231240 3943 231296
rect -960 231238 3943 231240
rect -960 231148 480 231238
rect 3877 231235 3943 231238
rect 38745 229938 38811 229941
rect 38745 229936 41124 229938
rect 38745 229880 38750 229936
rect 38806 229880 41124 229936
rect 38745 229878 41124 229880
rect 38745 229875 38811 229878
rect 544469 229802 544535 229805
rect 542892 229800 544535 229802
rect 542892 229744 544474 229800
rect 544530 229744 544535 229800
rect 542892 229742 544535 229744
rect 544469 229739 544535 229742
rect 580165 229122 580231 229125
rect 583520 229122 584960 229212
rect 580165 229120 584960 229122
rect 580165 229064 580170 229120
rect 580226 229064 584960 229120
rect 580165 229062 584960 229064
rect 580165 229059 580231 229062
rect 583520 228972 584960 229062
rect -960 226402 480 226492
rect 3141 226402 3207 226405
rect -960 226400 3207 226402
rect -960 226344 3146 226400
rect 3202 226344 3207 226400
rect -960 226342 3207 226344
rect -960 226252 480 226342
rect 3141 226339 3207 226342
rect 40309 225450 40375 225453
rect 40309 225448 41124 225450
rect 40309 225392 40314 225448
rect 40370 225392 41124 225448
rect 40309 225390 41124 225392
rect 40309 225387 40375 225390
rect 544745 225314 544811 225317
rect 542892 225312 544811 225314
rect 542892 225256 544750 225312
rect 544806 225256 544811 225312
rect 542892 225254 544811 225256
rect 544745 225251 544811 225254
rect 583520 224076 584960 224316
rect -960 221506 480 221596
rect 3877 221506 3943 221509
rect -960 221504 3943 221506
rect -960 221448 3882 221504
rect 3938 221448 3943 221504
rect -960 221446 3943 221448
rect -960 221356 480 221446
rect 3877 221443 3943 221446
rect 38837 220962 38903 220965
rect 38837 220960 41124 220962
rect 38837 220904 38842 220960
rect 38898 220904 41124 220960
rect 38837 220902 41124 220904
rect 38837 220899 38903 220902
rect 544745 220690 544811 220693
rect 542892 220688 544811 220690
rect 542892 220632 544750 220688
rect 544806 220632 544811 220688
rect 542892 220630 544811 220632
rect 544745 220627 544811 220630
rect 579797 219330 579863 219333
rect 583520 219330 584960 219420
rect 579797 219328 584960 219330
rect 579797 219272 579802 219328
rect 579858 219272 584960 219328
rect 579797 219270 584960 219272
rect 579797 219267 579863 219270
rect 583520 219180 584960 219270
rect -960 216610 480 216700
rect 3049 216610 3115 216613
rect -960 216608 3115 216610
rect -960 216552 3054 216608
rect 3110 216552 3115 216608
rect -960 216550 3115 216552
rect -960 216460 480 216550
rect 3049 216547 3115 216550
rect 40309 216338 40375 216341
rect 545573 216338 545639 216341
rect 40309 216336 41124 216338
rect 40309 216280 40314 216336
rect 40370 216280 41124 216336
rect 40309 216278 41124 216280
rect 542892 216336 545639 216338
rect 542892 216280 545578 216336
rect 545634 216280 545639 216336
rect 542892 216278 545639 216280
rect 40309 216275 40375 216278
rect 545573 216275 545639 216278
rect 580165 214162 580231 214165
rect 583520 214162 584960 214252
rect 580165 214160 584960 214162
rect 580165 214104 580170 214160
rect 580226 214104 584960 214160
rect 580165 214102 584960 214104
rect 580165 214099 580231 214102
rect 583520 214012 584960 214102
rect 40585 211986 40651 211989
rect 40585 211984 41124 211986
rect 40585 211928 40590 211984
rect 40646 211928 41124 211984
rect 40585 211926 41124 211928
rect 40585 211923 40651 211926
rect 544469 211714 544535 211717
rect 542892 211712 544535 211714
rect 542892 211656 544474 211712
rect 544530 211656 544535 211712
rect 542892 211654 544535 211656
rect 544469 211651 544535 211654
rect -960 211442 480 211532
rect 3601 211442 3667 211445
rect -960 211440 3667 211442
rect -960 211384 3606 211440
rect 3662 211384 3667 211440
rect -960 211382 3667 211384
rect -960 211292 480 211382
rect 3601 211379 3667 211382
rect 579981 209266 580047 209269
rect 583520 209266 584960 209356
rect 579981 209264 584960 209266
rect 579981 209208 579986 209264
rect 580042 209208 584960 209264
rect 579981 209206 584960 209208
rect 579981 209203 580047 209206
rect 583520 209116 584960 209206
rect 38837 207770 38903 207773
rect 38837 207768 41124 207770
rect 38837 207712 38842 207768
rect 38898 207712 41124 207768
rect 38837 207710 41124 207712
rect 38837 207707 38903 207710
rect 544745 207498 544811 207501
rect 542892 207496 544811 207498
rect 542892 207440 544750 207496
rect 544806 207440 544811 207496
rect 542892 207438 544811 207440
rect 544745 207435 544811 207438
rect -960 206546 480 206636
rect 3785 206546 3851 206549
rect -960 206544 3851 206546
rect -960 206488 3790 206544
rect 3846 206488 3851 206544
rect -960 206486 3851 206488
rect -960 206396 480 206486
rect 3785 206483 3851 206486
rect 580349 204370 580415 204373
rect 583520 204370 584960 204460
rect 580349 204368 584960 204370
rect 580349 204312 580354 204368
rect 580410 204312 584960 204368
rect 580349 204310 584960 204312
rect 580349 204307 580415 204310
rect 583520 204220 584960 204310
rect 39481 203146 39547 203149
rect 39481 203144 41124 203146
rect 39481 203088 39486 203144
rect 39542 203088 41124 203144
rect 39481 203086 41124 203088
rect 39481 203083 39547 203086
rect 542862 202194 542922 202708
rect 542997 202194 543063 202197
rect 542862 202192 543063 202194
rect 542862 202136 543002 202192
rect 543058 202136 543063 202192
rect 542862 202134 543063 202136
rect 542997 202131 543063 202134
rect -960 201650 480 201740
rect 3141 201650 3207 201653
rect -960 201648 3207 201650
rect -960 201592 3146 201648
rect 3202 201592 3207 201648
rect -960 201590 3207 201592
rect -960 201500 480 201590
rect 3141 201587 3207 201590
rect 580165 199474 580231 199477
rect 583520 199474 584960 199564
rect 580165 199472 584960 199474
rect 580165 199416 580170 199472
rect 580226 199416 584960 199472
rect 580165 199414 584960 199416
rect 580165 199411 580231 199414
rect 583520 199324 584960 199414
rect 39757 198794 39823 198797
rect 39757 198792 41124 198794
rect 39757 198736 39762 198792
rect 39818 198736 41124 198792
rect 39757 198734 41124 198736
rect 39757 198731 39823 198734
rect 543089 198386 543155 198389
rect 542892 198384 543155 198386
rect 542892 198328 543094 198384
rect 543150 198328 543155 198384
rect 542892 198326 543155 198328
rect 543089 198323 543155 198326
rect -960 196754 480 196844
rect 3141 196754 3207 196757
rect -960 196752 3207 196754
rect -960 196696 3146 196752
rect 3202 196696 3207 196752
rect -960 196694 3207 196696
rect -960 196604 480 196694
rect 3141 196691 3207 196694
rect 580165 194578 580231 194581
rect 583520 194578 584960 194668
rect 580165 194576 584960 194578
rect 580165 194520 580170 194576
rect 580226 194520 584960 194576
rect 580165 194518 584960 194520
rect 580165 194515 580231 194518
rect 583520 194428 584960 194518
rect 38837 194034 38903 194037
rect 38837 194032 41124 194034
rect 38837 193976 38842 194032
rect 38898 193976 41124 194032
rect 38837 193974 41124 193976
rect 38837 193971 38903 193974
rect 541942 193357 542002 193732
rect 541893 193352 542002 193357
rect 541893 193296 541898 193352
rect 541954 193296 542002 193352
rect 541893 193294 542002 193296
rect 541893 193291 541959 193294
rect -960 191858 480 191948
rect 3877 191858 3943 191861
rect -960 191856 3943 191858
rect -960 191800 3882 191856
rect 3938 191800 3943 191856
rect -960 191798 3943 191800
rect -960 191708 480 191798
rect 3877 191795 3943 191798
rect 543590 191660 543596 191724
rect 543660 191722 543666 191724
rect 544469 191722 544535 191725
rect 543660 191720 544535 191722
rect 543660 191664 544474 191720
rect 544530 191664 544535 191720
rect 543660 191662 544535 191664
rect 543660 191660 543666 191662
rect 544469 191659 544535 191662
rect 39481 189818 39547 189821
rect 39481 189816 41124 189818
rect 39481 189760 39486 189816
rect 39542 189760 41124 189816
rect 39481 189758 41124 189760
rect 39481 189755 39547 189758
rect 579613 189682 579679 189685
rect 583520 189682 584960 189772
rect 579613 189680 584960 189682
rect 579613 189624 579618 189680
rect 579674 189624 584960 189680
rect 579613 189622 584960 189624
rect 579613 189619 579679 189622
rect 583520 189532 584960 189622
rect 545665 189410 545731 189413
rect 542892 189408 545731 189410
rect 542892 189352 545670 189408
rect 545726 189352 545731 189408
rect 542892 189350 545731 189352
rect 545665 189347 545731 189350
rect -960 186962 480 187052
rect 3141 186962 3207 186965
rect -960 186960 3207 186962
rect -960 186904 3146 186960
rect 3202 186904 3207 186960
rect -960 186902 3207 186904
rect -960 186812 480 186902
rect 3141 186899 3207 186902
rect 38837 185058 38903 185061
rect 38837 185056 41124 185058
rect 38837 185000 38842 185056
rect 38898 185000 41124 185056
rect 38837 184998 41124 185000
rect 38837 184995 38903 184998
rect 544745 184786 544811 184789
rect 542892 184784 544811 184786
rect 542892 184728 544750 184784
rect 544806 184728 544811 184784
rect 542892 184726 544811 184728
rect 544745 184723 544811 184726
rect 580165 184786 580231 184789
rect 583520 184786 584960 184876
rect 580165 184784 584960 184786
rect 580165 184728 580170 184784
rect 580226 184728 584960 184784
rect 580165 184726 584960 184728
rect 580165 184723 580231 184726
rect 583520 184636 584960 184726
rect -960 182066 480 182156
rect 3141 182066 3207 182069
rect -960 182064 3207 182066
rect -960 182008 3146 182064
rect 3202 182008 3207 182064
rect -960 182006 3207 182008
rect -960 181916 480 182006
rect 3141 182003 3207 182006
rect 39113 180842 39179 180845
rect 39113 180840 41124 180842
rect 39113 180784 39118 180840
rect 39174 180784 41124 180840
rect 39113 180782 41124 180784
rect 39113 180779 39179 180782
rect 543825 180570 543891 180573
rect 542892 180568 543891 180570
rect 542892 180512 543830 180568
rect 543886 180512 543891 180568
rect 542892 180510 543891 180512
rect 543825 180507 543891 180510
rect 579981 179890 580047 179893
rect 583520 179890 584960 179980
rect 579981 179888 584960 179890
rect 579981 179832 579986 179888
rect 580042 179832 584960 179888
rect 579981 179830 584960 179832
rect 579981 179827 580047 179830
rect 583520 179740 584960 179830
rect -960 177170 480 177260
rect 3049 177170 3115 177173
rect -960 177168 3115 177170
rect -960 177112 3054 177168
rect 3110 177112 3115 177168
rect -960 177110 3115 177112
rect -960 177020 480 177110
rect 3049 177107 3115 177110
rect 38837 176218 38903 176221
rect 38837 176216 41124 176218
rect 38837 176160 38842 176216
rect 38898 176160 41124 176216
rect 38837 176158 41124 176160
rect 38837 176155 38903 176158
rect 544745 175946 544811 175949
rect 542892 175944 544811 175946
rect 542892 175888 544750 175944
rect 544806 175888 544811 175944
rect 542892 175886 544811 175888
rect 544745 175883 544811 175886
rect 579613 174994 579679 174997
rect 583520 174994 584960 175084
rect 579613 174992 584960 174994
rect 579613 174936 579618 174992
rect 579674 174936 584960 174992
rect 579613 174934 584960 174936
rect 579613 174931 579679 174934
rect 583520 174844 584960 174934
rect -960 172274 480 172364
rect 3049 172274 3115 172277
rect -960 172272 3115 172274
rect -960 172216 3054 172272
rect 3110 172216 3115 172272
rect -960 172214 3115 172216
rect -960 172124 480 172214
rect 3049 172211 3115 172214
rect 39481 171730 39547 171733
rect 39481 171728 41124 171730
rect 39481 171672 39486 171728
rect 39542 171672 41124 171728
rect 39481 171670 41124 171672
rect 39481 171667 39547 171670
rect 544469 171458 544535 171461
rect 542892 171456 544535 171458
rect 542892 171400 544474 171456
rect 544530 171400 544535 171456
rect 542892 171398 544535 171400
rect 544469 171395 544535 171398
rect 580901 170098 580967 170101
rect 583520 170098 584960 170188
rect 580901 170096 584960 170098
rect 580901 170040 580906 170096
rect 580962 170040 584960 170096
rect 580901 170038 584960 170040
rect 580901 170035 580967 170038
rect 583520 169948 584960 170038
rect -960 167378 480 167468
rect 3141 167378 3207 167381
rect -960 167376 3207 167378
rect -960 167320 3146 167376
rect 3202 167320 3207 167376
rect -960 167318 3207 167320
rect -960 167228 480 167318
rect 3141 167315 3207 167318
rect 38837 167242 38903 167245
rect 543825 167242 543891 167245
rect 38837 167240 41124 167242
rect 38837 167184 38842 167240
rect 38898 167184 41124 167240
rect 38837 167182 41124 167184
rect 542892 167240 543891 167242
rect 542892 167184 543830 167240
rect 543886 167184 543891 167240
rect 542892 167182 543891 167184
rect 38837 167179 38903 167182
rect 543825 167179 543891 167182
rect 579981 165202 580047 165205
rect 583520 165202 584960 165292
rect 579981 165200 584960 165202
rect 579981 165144 579986 165200
rect 580042 165144 584960 165200
rect 579981 165142 584960 165144
rect 579981 165139 580047 165142
rect 583520 165052 584960 165142
rect 38837 162754 38903 162757
rect 38837 162752 41124 162754
rect 38837 162696 38842 162752
rect 38898 162696 41124 162752
rect 38837 162694 41124 162696
rect 38837 162691 38903 162694
rect -960 162482 480 162572
rect 2773 162482 2839 162485
rect 543825 162482 543891 162485
rect -960 162480 2839 162482
rect -960 162424 2778 162480
rect 2834 162424 2839 162480
rect -960 162422 2839 162424
rect 542892 162480 543891 162482
rect 542892 162424 543830 162480
rect 543886 162424 543891 162480
rect 542892 162422 543891 162424
rect -960 162332 480 162422
rect 2773 162419 2839 162422
rect 543825 162419 543891 162422
rect 580165 160034 580231 160037
rect 583520 160034 584960 160124
rect 580165 160032 584960 160034
rect 580165 159976 580170 160032
rect 580226 159976 584960 160032
rect 580165 159974 584960 159976
rect 580165 159971 580231 159974
rect 583520 159884 584960 159974
rect 544745 158266 544811 158269
rect 542892 158264 544811 158266
rect 542892 158208 544750 158264
rect 544806 158208 544811 158264
rect 542892 158206 544811 158208
rect 544745 158203 544811 158206
rect 39297 158130 39363 158133
rect 39297 158128 41124 158130
rect 39297 158072 39302 158128
rect 39358 158072 41124 158128
rect 39297 158070 41124 158072
rect 39297 158067 39363 158070
rect -960 157314 480 157404
rect 3417 157314 3483 157317
rect -960 157312 3483 157314
rect -960 157256 3422 157312
rect 3478 157256 3483 157312
rect -960 157254 3483 157256
rect -960 157164 480 157254
rect 3417 157251 3483 157254
rect 579613 155138 579679 155141
rect 583520 155138 584960 155228
rect 579613 155136 584960 155138
rect 579613 155080 579618 155136
rect 579674 155080 584960 155136
rect 579613 155078 584960 155080
rect 579613 155075 579679 155078
rect 583520 154988 584960 155078
rect 39941 153778 40007 153781
rect 39941 153776 41124 153778
rect 39941 153720 39946 153776
rect 40002 153720 41124 153776
rect 39941 153718 41124 153720
rect 39941 153715 40007 153718
rect 543273 153506 543339 153509
rect 542892 153504 543339 153506
rect 542892 153448 543278 153504
rect 543334 153448 543339 153504
rect 542892 153446 543339 153448
rect 543273 153443 543339 153446
rect -960 152268 480 152508
rect 541750 150452 541756 150516
rect 541820 150514 541826 150516
rect 543825 150514 543891 150517
rect 541820 150512 543891 150514
rect 541820 150456 543830 150512
rect 543886 150456 543891 150512
rect 541820 150454 543891 150456
rect 541820 150452 541826 150454
rect 543825 150451 543891 150454
rect 579613 150242 579679 150245
rect 583520 150242 584960 150332
rect 579613 150240 584960 150242
rect 579613 150184 579618 150240
rect 579674 150184 584960 150240
rect 579613 150182 584960 150184
rect 579613 150179 579679 150182
rect 583520 150092 584960 150182
rect 40033 149562 40099 149565
rect 40033 149560 41124 149562
rect 40033 149504 40038 149560
rect 40094 149504 41124 149560
rect 40033 149502 41124 149504
rect 40033 149499 40099 149502
rect 544653 149290 544719 149293
rect 542892 149288 544719 149290
rect 542892 149232 544658 149288
rect 544714 149232 544719 149288
rect 542892 149230 544719 149232
rect 544653 149227 544719 149230
rect -960 147522 480 147612
rect 3417 147522 3483 147525
rect -960 147520 3483 147522
rect -960 147464 3422 147520
rect 3478 147464 3483 147520
rect -960 147462 3483 147464
rect -960 147372 480 147462
rect 3417 147459 3483 147462
rect 583520 145196 584960 145436
rect 39205 144802 39271 144805
rect 39205 144800 41124 144802
rect 39205 144744 39210 144800
rect 39266 144744 41124 144800
rect 39205 144742 41124 144744
rect 39205 144739 39271 144742
rect 541942 143989 542002 144500
rect 541942 143984 542051 143989
rect 541942 143928 541990 143984
rect 542046 143928 542051 143984
rect 541942 143926 542051 143928
rect 541985 143923 542051 143926
rect -960 142626 480 142716
rect 2773 142626 2839 142629
rect -960 142624 2839 142626
rect -960 142568 2778 142624
rect 2834 142568 2839 142624
rect -960 142566 2839 142568
rect -960 142476 480 142566
rect 2773 142563 2839 142566
rect 38929 140450 38995 140453
rect 580165 140450 580231 140453
rect 583520 140450 584960 140540
rect 38929 140448 41124 140450
rect 38929 140392 38934 140448
rect 38990 140392 41124 140448
rect 38929 140390 41124 140392
rect 580165 140448 584960 140450
rect 580165 140392 580170 140448
rect 580226 140392 584960 140448
rect 580165 140390 584960 140392
rect 38929 140387 38995 140390
rect 580165 140387 580231 140390
rect 583520 140300 584960 140390
rect 543181 140178 543247 140181
rect 542892 140176 543247 140178
rect 542892 140120 543186 140176
rect 543242 140120 543247 140176
rect 542892 140118 543247 140120
rect 543181 140115 543247 140118
rect 542854 139436 542860 139500
rect 542924 139498 542930 139500
rect 543825 139498 543891 139501
rect 542924 139496 543891 139498
rect 542924 139440 543830 139496
rect 543886 139440 543891 139496
rect 542924 139438 543891 139440
rect 542924 139436 542930 139438
rect 543825 139435 543891 139438
rect -960 137730 480 137820
rect 3417 137730 3483 137733
rect -960 137728 3483 137730
rect -960 137672 3422 137728
rect 3478 137672 3483 137728
rect -960 137670 3483 137672
rect -960 137580 480 137670
rect 3417 137667 3483 137670
rect 39389 135826 39455 135829
rect 39389 135824 41124 135826
rect 39389 135768 39394 135824
rect 39450 135768 41124 135824
rect 39389 135766 41124 135768
rect 39389 135763 39455 135766
rect 544326 135554 544332 135556
rect 542892 135494 544332 135554
rect 544326 135492 544332 135494
rect 544396 135492 544402 135556
rect 579613 135554 579679 135557
rect 583520 135554 584960 135644
rect 579613 135552 584960 135554
rect 579613 135496 579618 135552
rect 579674 135496 584960 135552
rect 579613 135494 584960 135496
rect 579613 135491 579679 135494
rect 583520 135404 584960 135494
rect -960 132834 480 132924
rect 3417 132834 3483 132837
rect -960 132832 3483 132834
rect -960 132776 3422 132832
rect 3478 132776 3483 132832
rect -960 132774 3483 132776
rect -960 132684 480 132774
rect 3417 132771 3483 132774
rect 38837 131610 38903 131613
rect 38837 131608 41124 131610
rect 38837 131552 38842 131608
rect 38898 131552 41124 131608
rect 38837 131550 41124 131552
rect 38837 131547 38903 131550
rect 543825 131338 543891 131341
rect 542892 131336 543891 131338
rect 542892 131280 543830 131336
rect 543886 131280 543891 131336
rect 542892 131278 543891 131280
rect 543825 131275 543891 131278
rect 579797 130658 579863 130661
rect 583520 130658 584960 130748
rect 579797 130656 584960 130658
rect 579797 130600 579802 130656
rect 579858 130600 584960 130656
rect 579797 130598 584960 130600
rect 579797 130595 579863 130598
rect 583520 130508 584960 130598
rect -960 127938 480 128028
rect 3233 127938 3299 127941
rect -960 127936 3299 127938
rect -960 127880 3238 127936
rect 3294 127880 3299 127936
rect -960 127878 3299 127880
rect -960 127788 480 127878
rect 3233 127875 3299 127878
rect 40033 126850 40099 126853
rect 40033 126848 41124 126850
rect 40033 126792 40038 126848
rect 40094 126792 41124 126848
rect 40033 126790 41124 126792
rect 40033 126787 40099 126790
rect 545021 126578 545087 126581
rect 542892 126576 545087 126578
rect 542892 126520 545026 126576
rect 545082 126520 545087 126576
rect 542892 126518 545087 126520
rect 545021 126515 545087 126518
rect 580717 125762 580783 125765
rect 583520 125762 584960 125852
rect 580717 125760 584960 125762
rect 580717 125704 580722 125760
rect 580778 125704 584960 125760
rect 580717 125702 584960 125704
rect 580717 125699 580783 125702
rect 583520 125612 584960 125702
rect -960 123042 480 123132
rect 3601 123042 3667 123045
rect -960 123040 3667 123042
rect -960 122984 3606 123040
rect 3662 122984 3667 123040
rect -960 122982 3667 122984
rect -960 122892 480 122982
rect 3601 122979 3667 122982
rect 38101 122634 38167 122637
rect 38101 122632 41124 122634
rect 38101 122576 38106 122632
rect 38162 122576 41124 122632
rect 38101 122574 41124 122576
rect 38101 122571 38167 122574
rect 544469 122226 544535 122229
rect 542892 122224 544535 122226
rect 542892 122168 544474 122224
rect 544530 122168 544535 122224
rect 542892 122166 544535 122168
rect 544469 122163 544535 122166
rect 580165 120866 580231 120869
rect 583520 120866 584960 120956
rect 580165 120864 584960 120866
rect 580165 120808 580170 120864
rect 580226 120808 584960 120864
rect 580165 120806 584960 120808
rect 580165 120803 580231 120806
rect 583520 120716 584960 120806
rect -960 118146 480 118236
rect 3601 118146 3667 118149
rect -960 118144 3667 118146
rect -960 118088 3606 118144
rect 3662 118088 3667 118144
rect -960 118086 3667 118088
rect -960 117996 480 118086
rect 3601 118083 3667 118086
rect 39614 117948 39620 118012
rect 39684 118010 39690 118012
rect 39684 117950 41124 118010
rect 39684 117948 39690 117950
rect 542126 117333 542186 117572
rect 542126 117328 542235 117333
rect 542126 117272 542174 117328
rect 542230 117272 542235 117328
rect 542126 117270 542235 117272
rect 542169 117267 542235 117270
rect 579613 115970 579679 115973
rect 583520 115970 584960 116060
rect 579613 115968 584960 115970
rect 579613 115912 579618 115968
rect 579674 115912 584960 115968
rect 579613 115910 584960 115912
rect 579613 115907 579679 115910
rect 583520 115820 584960 115910
rect 38837 113658 38903 113661
rect 38837 113656 41124 113658
rect 38837 113600 38842 113656
rect 38898 113600 41124 113656
rect 38837 113598 41124 113600
rect 38837 113595 38903 113598
rect 544653 113386 544719 113389
rect 542892 113384 544719 113386
rect -960 113250 480 113340
rect 542892 113328 544658 113384
rect 544714 113328 544719 113384
rect 542892 113326 544719 113328
rect 544653 113323 544719 113326
rect 3049 113250 3115 113253
rect -960 113248 3115 113250
rect -960 113192 3054 113248
rect 3110 113192 3115 113248
rect -960 113190 3115 113192
rect -960 113100 480 113190
rect 3049 113187 3115 113190
rect 580165 111074 580231 111077
rect 583520 111074 584960 111164
rect 580165 111072 584960 111074
rect 580165 111016 580170 111072
rect 580226 111016 584960 111072
rect 580165 111014 584960 111016
rect 580165 111011 580231 111014
rect 583520 110924 584960 111014
rect 38837 109034 38903 109037
rect 543733 109034 543799 109037
rect 38837 109032 41124 109034
rect 38837 108976 38842 109032
rect 38898 108976 41124 109032
rect 38837 108974 41124 108976
rect 542892 109032 543799 109034
rect 542892 108976 543738 109032
rect 543794 108976 543799 109032
rect 542892 108974 543799 108976
rect 38837 108971 38903 108974
rect 543733 108971 543799 108974
rect -960 108354 480 108444
rect 3141 108354 3207 108357
rect -960 108352 3207 108354
rect -960 108296 3146 108352
rect 3202 108296 3207 108352
rect -960 108294 3207 108296
rect -960 108204 480 108294
rect 3141 108291 3207 108294
rect 580165 105906 580231 105909
rect 583520 105906 584960 105996
rect 580165 105904 584960 105906
rect 580165 105848 580170 105904
rect 580226 105848 584960 105904
rect 580165 105846 584960 105848
rect 580165 105843 580231 105846
rect 583520 105756 584960 105846
rect 39849 104546 39915 104549
rect 39849 104544 41124 104546
rect 39849 104488 39854 104544
rect 39910 104488 41124 104544
rect 39849 104486 41124 104488
rect 39849 104483 39915 104486
rect 543733 104274 543799 104277
rect 542892 104272 543799 104274
rect 542892 104216 543738 104272
rect 543794 104216 543799 104272
rect 542892 104214 543799 104216
rect 543733 104211 543799 104214
rect -960 103186 480 103276
rect 3325 103186 3391 103189
rect -960 103184 3391 103186
rect -960 103128 3330 103184
rect 3386 103128 3391 103184
rect -960 103126 3391 103128
rect -960 103036 480 103126
rect 3325 103123 3391 103126
rect 579613 101010 579679 101013
rect 583520 101010 584960 101100
rect 579613 101008 584960 101010
rect 579613 100952 579618 101008
rect 579674 100952 584960 101008
rect 579613 100950 584960 100952
rect 579613 100947 579679 100950
rect 583520 100860 584960 100950
rect 39941 99922 40007 99925
rect 544653 99922 544719 99925
rect 39941 99920 41124 99922
rect 39941 99864 39946 99920
rect 40002 99864 41124 99920
rect 39941 99862 41124 99864
rect 542892 99920 544719 99922
rect 542892 99864 544658 99920
rect 544714 99864 544719 99920
rect 542892 99862 544719 99864
rect 39941 99859 40007 99862
rect 544653 99859 544719 99862
rect -960 98140 480 98380
rect 578969 96114 579035 96117
rect 583520 96114 584960 96204
rect 578969 96112 584960 96114
rect 578969 96056 578974 96112
rect 579030 96056 584960 96112
rect 578969 96054 584960 96056
rect 578969 96051 579035 96054
rect 583520 95964 584960 96054
rect 39021 95570 39087 95573
rect 39021 95568 41124 95570
rect 39021 95512 39026 95568
rect 39082 95512 41124 95568
rect 39021 95510 41124 95512
rect 39021 95507 39087 95510
rect 542126 95165 542186 95268
rect 542077 95160 542186 95165
rect 542077 95104 542082 95160
rect 542138 95104 542186 95160
rect 542077 95102 542186 95104
rect 542077 95099 542143 95102
rect -960 93394 480 93484
rect 2773 93394 2839 93397
rect -960 93392 2839 93394
rect -960 93336 2778 93392
rect 2834 93336 2839 93392
rect -960 93334 2839 93336
rect -960 93244 480 93334
rect 2773 93331 2839 93334
rect 38929 91218 38995 91221
rect 38929 91216 41124 91218
rect 38929 91160 38934 91216
rect 38990 91160 41124 91216
rect 38929 91158 41124 91160
rect 38929 91155 38995 91158
rect 583520 91068 584960 91308
rect 544745 90946 544811 90949
rect 542892 90944 544811 90946
rect 542892 90888 544750 90944
rect 544806 90888 544811 90944
rect 542892 90886 544811 90888
rect 544745 90883 544811 90886
rect -960 88498 480 88588
rect 3601 88498 3667 88501
rect -960 88496 3667 88498
rect -960 88440 3606 88496
rect 3662 88440 3667 88496
rect -960 88438 3667 88440
rect -960 88348 480 88438
rect 3601 88435 3667 88438
rect 38837 86594 38903 86597
rect 38837 86592 41124 86594
rect 38837 86536 38842 86592
rect 38898 86536 41124 86592
rect 38837 86534 41124 86536
rect 38837 86531 38903 86534
rect 543457 86322 543523 86325
rect 542892 86320 543523 86322
rect 542892 86264 543462 86320
rect 543518 86264 543523 86320
rect 542892 86262 543523 86264
rect 543457 86259 543523 86262
rect 578877 86322 578943 86325
rect 583520 86322 584960 86412
rect 578877 86320 584960 86322
rect 578877 86264 578882 86320
rect 578938 86264 584960 86320
rect 578877 86262 584960 86264
rect 578877 86259 578943 86262
rect 583520 86172 584960 86262
rect -960 83602 480 83692
rect 3325 83602 3391 83605
rect -960 83600 3391 83602
rect -960 83544 3330 83600
rect 3386 83544 3391 83600
rect -960 83542 3391 83544
rect -960 83452 480 83542
rect 3325 83539 3391 83542
rect 39113 82242 39179 82245
rect 39113 82240 41124 82242
rect 39113 82184 39118 82240
rect 39174 82184 41124 82240
rect 39113 82182 41124 82184
rect 39113 82179 39179 82182
rect 543825 81970 543891 81973
rect 542892 81968 543891 81970
rect 542892 81912 543830 81968
rect 543886 81912 543891 81968
rect 542892 81910 543891 81912
rect 543825 81907 543891 81910
rect 580165 81426 580231 81429
rect 583520 81426 584960 81516
rect 580165 81424 584960 81426
rect 580165 81368 580170 81424
rect 580226 81368 584960 81424
rect 580165 81366 584960 81368
rect 580165 81363 580231 81366
rect 583520 81276 584960 81366
rect -960 78706 480 78796
rect 2773 78706 2839 78709
rect -960 78704 2839 78706
rect -960 78648 2778 78704
rect 2834 78648 2839 78704
rect -960 78646 2839 78648
rect -960 78556 480 78646
rect 2773 78643 2839 78646
rect 40033 77618 40099 77621
rect 40033 77616 41124 77618
rect 40033 77560 40038 77616
rect 40094 77560 41124 77616
rect 40033 77558 41124 77560
rect 40033 77555 40099 77558
rect 543733 77346 543799 77349
rect 542892 77344 543799 77346
rect 542892 77288 543738 77344
rect 543794 77288 543799 77344
rect 542892 77286 543799 77288
rect 543733 77283 543799 77286
rect 583520 76380 584960 76620
rect -960 73810 480 73900
rect 3325 73810 3391 73813
rect -960 73808 3391 73810
rect -960 73752 3330 73808
rect 3386 73752 3391 73808
rect -960 73750 3391 73752
rect -960 73660 480 73750
rect 3325 73747 3391 73750
rect 39849 73266 39915 73269
rect 39849 73264 41124 73266
rect 39849 73208 39854 73264
rect 39910 73208 41124 73264
rect 39849 73206 41124 73208
rect 39849 73203 39915 73206
rect 545665 72994 545731 72997
rect 542892 72992 545731 72994
rect 542892 72936 545670 72992
rect 545726 72936 545731 72992
rect 542892 72934 545731 72936
rect 545665 72931 545731 72934
rect 580809 71634 580875 71637
rect 583520 71634 584960 71724
rect 580809 71632 584960 71634
rect 580809 71576 580814 71632
rect 580870 71576 584960 71632
rect 580809 71574 584960 71576
rect 580809 71571 580875 71574
rect 583520 71484 584960 71574
rect -960 68914 480 69004
rect 3325 68914 3391 68917
rect -960 68912 3391 68914
rect -960 68856 3330 68912
rect 3386 68856 3391 68912
rect -960 68854 3391 68856
rect -960 68764 480 68854
rect 3325 68851 3391 68854
rect 38193 68778 38259 68781
rect 38193 68776 41124 68778
rect 38193 68720 38198 68776
rect 38254 68720 41124 68776
rect 38193 68718 41124 68720
rect 38193 68715 38259 68718
rect 543825 68506 543891 68509
rect 542892 68504 543891 68506
rect 542892 68448 543830 68504
rect 543886 68448 543891 68504
rect 542892 68446 543891 68448
rect 543825 68443 543891 68446
rect 580901 66738 580967 66741
rect 583520 66738 584960 66828
rect 580901 66736 584960 66738
rect 580901 66680 580906 66736
rect 580962 66680 584960 66736
rect 580901 66678 584960 66680
rect 580901 66675 580967 66678
rect 583520 66588 584960 66678
rect 39941 64290 40007 64293
rect 39941 64288 41124 64290
rect 39941 64232 39946 64288
rect 40002 64232 41124 64288
rect 39941 64230 41124 64232
rect 39941 64227 40007 64230
rect 543825 64154 543891 64157
rect 542892 64152 543891 64154
rect -960 64018 480 64108
rect 542892 64096 543830 64152
rect 543886 64096 543891 64152
rect 542892 64094 543891 64096
rect 543825 64091 543891 64094
rect 2773 64018 2839 64021
rect -960 64016 2839 64018
rect -960 63960 2778 64016
rect 2834 63960 2839 64016
rect -960 63958 2839 63960
rect -960 63868 480 63958
rect 2773 63955 2839 63958
rect 580165 61842 580231 61845
rect 583520 61842 584960 61932
rect 580165 61840 584960 61842
rect 580165 61784 580170 61840
rect 580226 61784 584960 61840
rect 580165 61782 584960 61784
rect 580165 61779 580231 61782
rect 583520 61692 584960 61782
rect 38837 59666 38903 59669
rect 38837 59664 41124 59666
rect 38837 59608 38842 59664
rect 38898 59608 41124 59664
rect 38837 59606 41124 59608
rect 38837 59603 38903 59606
rect 543825 59530 543891 59533
rect 542892 59528 543891 59530
rect 542892 59472 543830 59528
rect 543886 59472 543891 59528
rect 542892 59470 543891 59472
rect 543825 59467 543891 59470
rect -960 59122 480 59212
rect 3785 59122 3851 59125
rect -960 59120 3851 59122
rect -960 59064 3790 59120
rect 3846 59064 3851 59120
rect -960 59062 3851 59064
rect -960 58972 480 59062
rect 3785 59059 3851 59062
rect 580073 56946 580139 56949
rect 583520 56946 584960 57036
rect 580073 56944 584960 56946
rect 580073 56888 580078 56944
rect 580134 56888 584960 56944
rect 580073 56886 584960 56888
rect 580073 56883 580139 56886
rect 583520 56796 584960 56886
rect 39982 55388 39988 55452
rect 40052 55450 40058 55452
rect 40052 55390 41124 55450
rect 40052 55388 40058 55390
rect 543825 55042 543891 55045
rect 542892 55040 543891 55042
rect 542892 54984 543830 55040
rect 543886 54984 543891 55040
rect 542892 54982 543891 54984
rect 543825 54979 543891 54982
rect -960 54226 480 54316
rect 3325 54226 3391 54229
rect -960 54224 3391 54226
rect -960 54168 3330 54224
rect 3386 54168 3391 54224
rect -960 54166 3391 54168
rect -960 54076 480 54166
rect 3325 54163 3391 54166
rect 579981 51778 580047 51781
rect 583520 51778 584960 51868
rect 579981 51776 584960 51778
rect 579981 51720 579986 51776
rect 580042 51720 584960 51776
rect 579981 51718 584960 51720
rect 579981 51715 580047 51718
rect 583520 51628 584960 51718
rect 543825 50690 543891 50693
rect 542892 50688 543891 50690
rect 40953 50146 41019 50149
rect 41094 50146 41154 50660
rect 542892 50632 543830 50688
rect 543886 50632 543891 50688
rect 542892 50630 543891 50632
rect 543825 50627 543891 50630
rect 40953 50144 41154 50146
rect 40953 50088 40958 50144
rect 41014 50088 41154 50144
rect 40953 50086 41154 50088
rect 40953 50083 41019 50086
rect 541934 49540 541940 49604
rect 542004 49602 542010 49604
rect 544326 49602 544332 49604
rect 542004 49542 544332 49602
rect 542004 49540 542010 49542
rect 544326 49540 544332 49542
rect 544396 49540 544402 49604
rect -960 49058 480 49148
rect 2773 49058 2839 49061
rect -960 49056 2839 49058
rect -960 49000 2778 49056
rect 2834 49000 2839 49056
rect -960 48998 2839 49000
rect -960 48908 480 48998
rect 2773 48995 2839 48998
rect 579981 46882 580047 46885
rect 583520 46882 584960 46972
rect 579981 46880 584960 46882
rect 579981 46824 579986 46880
rect 580042 46824 584960 46880
rect 579981 46822 584960 46824
rect 579981 46819 580047 46822
rect 583520 46732 584960 46822
rect 41094 45658 41154 46308
rect 544653 46202 544719 46205
rect 542892 46200 544719 46202
rect 542892 46144 544658 46200
rect 544714 46144 544719 46200
rect 542892 46142 544719 46144
rect 544653 46139 544719 46142
rect 40542 45598 41154 45658
rect 40542 45525 40602 45598
rect 40493 45520 40602 45525
rect 40493 45464 40498 45520
rect 40554 45464 40602 45520
rect 40493 45462 40602 45464
rect 40493 45459 40559 45462
rect 40166 44644 40172 44708
rect 40236 44706 40242 44708
rect 580717 44706 580783 44709
rect 40236 44704 580783 44706
rect 40236 44648 580722 44704
rect 580778 44648 580783 44704
rect 40236 44646 580783 44648
rect 40236 44644 40242 44646
rect 580717 44643 580783 44646
rect 10961 44570 11027 44573
rect 542670 44570 542676 44572
rect 10961 44568 542676 44570
rect 10961 44512 10966 44568
rect 11022 44512 542676 44568
rect 10961 44510 542676 44512
rect 10961 44507 11027 44510
rect 542670 44508 542676 44510
rect 542740 44508 542746 44572
rect 38101 44434 38167 44437
rect 541750 44434 541756 44436
rect 38101 44432 541756 44434
rect 38101 44376 38106 44432
rect 38162 44376 541756 44432
rect 38101 44374 541756 44376
rect 38101 44371 38167 44374
rect 541750 44372 541756 44374
rect 541820 44372 541826 44436
rect 41873 44298 41939 44301
rect 541566 44298 541572 44300
rect 41873 44296 541572 44298
rect -960 44162 480 44252
rect 41873 44240 41878 44296
rect 41934 44240 541572 44296
rect 41873 44238 541572 44240
rect 41873 44235 41939 44238
rect 541566 44236 541572 44238
rect 541636 44236 541642 44300
rect 4061 44162 4127 44165
rect -960 44160 4127 44162
rect -960 44104 4066 44160
rect 4122 44104 4127 44160
rect -960 44102 4127 44104
rect -960 44012 480 44102
rect 4061 44099 4127 44102
rect 38878 44100 38884 44164
rect 38948 44162 38954 44164
rect 552013 44162 552079 44165
rect 38948 44160 552079 44162
rect 38948 44104 552018 44160
rect 552074 44104 552079 44160
rect 38948 44102 552079 44104
rect 38948 44100 38954 44102
rect 552013 44099 552079 44102
rect 38837 44026 38903 44029
rect 541934 44026 541940 44028
rect 38837 44024 541940 44026
rect 38837 43968 38842 44024
rect 38898 43968 541940 44024
rect 38837 43966 541940 43968
rect 38837 43963 38903 43966
rect 541934 43964 541940 43966
rect 542004 43964 542010 44028
rect 55990 43828 55996 43892
rect 56060 43890 56066 43892
rect 122598 43890 122604 43892
rect 56060 43830 122604 43890
rect 56060 43828 56066 43830
rect 122598 43828 122604 43830
rect 122668 43828 122674 43892
rect 283966 43828 283972 43892
rect 284036 43890 284042 43892
rect 354806 43890 354812 43892
rect 284036 43830 354812 43890
rect 284036 43828 284042 43830
rect 354806 43828 354812 43830
rect 354876 43828 354882 43892
rect 53230 43692 53236 43756
rect 53300 43754 53306 43756
rect 207606 43754 207612 43756
rect 53300 43694 207612 43754
rect 53300 43692 53306 43694
rect 207606 43692 207612 43694
rect 207676 43692 207682 43756
rect 223982 43692 223988 43756
rect 224052 43754 224058 43756
rect 351862 43754 351868 43756
rect 224052 43694 351868 43754
rect 224052 43692 224058 43694
rect 351862 43692 351868 43694
rect 351932 43692 351938 43756
rect 39430 43556 39436 43620
rect 39500 43618 39506 43620
rect 554773 43618 554839 43621
rect 39500 43616 554839 43618
rect 39500 43560 554778 43616
rect 554834 43560 554839 43616
rect 39500 43558 554839 43560
rect 39500 43556 39506 43558
rect 554773 43555 554839 43558
rect 3877 43482 3943 43485
rect 544142 43482 544148 43484
rect 3877 43480 544148 43482
rect 3877 43424 3882 43480
rect 3938 43424 544148 43480
rect 3877 43422 544148 43424
rect 3877 43419 3943 43422
rect 544142 43420 544148 43422
rect 544212 43420 544218 43484
rect 295926 43284 295932 43348
rect 295996 43346 296002 43348
rect 355174 43346 355180 43348
rect 295996 43286 355180 43346
rect 295996 43284 296002 43286
rect 355174 43284 355180 43286
rect 355244 43284 355250 43348
rect 313222 43148 313228 43212
rect 313292 43210 313298 43212
rect 352414 43210 352420 43212
rect 313292 43150 352420 43210
rect 313292 43148 313298 43150
rect 352414 43148 352420 43150
rect 352484 43148 352490 43212
rect 54886 42332 54892 42396
rect 54956 42394 54962 42396
rect 59261 42394 59327 42397
rect 223941 42396 224007 42397
rect 284017 42396 284083 42397
rect 223941 42394 223988 42396
rect 54956 42392 59327 42394
rect 54956 42336 59266 42392
rect 59322 42336 59327 42392
rect 54956 42334 59327 42336
rect 223896 42392 223988 42394
rect 223896 42336 223946 42392
rect 223896 42334 223988 42336
rect 54956 42332 54962 42334
rect 59261 42331 59327 42334
rect 223941 42332 223988 42334
rect 224052 42332 224058 42396
rect 283966 42332 283972 42396
rect 284036 42394 284083 42396
rect 284036 42392 284128 42394
rect 284078 42336 284128 42392
rect 284036 42334 284128 42336
rect 284036 42332 284083 42334
rect 370446 42332 370452 42396
rect 370516 42394 370522 42396
rect 371693 42394 371759 42397
rect 405549 42396 405615 42397
rect 405549 42394 405596 42396
rect 370516 42392 371759 42394
rect 370516 42336 371698 42392
rect 371754 42336 371759 42392
rect 370516 42334 371759 42336
rect 405504 42392 405596 42394
rect 405504 42336 405554 42392
rect 405504 42334 405596 42336
rect 370516 42332 370522 42334
rect 223941 42331 224007 42332
rect 284017 42331 284083 42332
rect 371693 42331 371759 42334
rect 405549 42332 405596 42334
rect 405660 42332 405666 42396
rect 405549 42331 405615 42332
rect 54702 42196 54708 42260
rect 54772 42258 54778 42260
rect 68001 42258 68067 42261
rect 54772 42256 68067 42258
rect 54772 42200 68006 42256
rect 68062 42200 68067 42256
rect 54772 42198 68067 42200
rect 54772 42196 54778 42198
rect 68001 42195 68067 42198
rect 53414 42060 53420 42124
rect 53484 42122 53490 42124
rect 157425 42122 157491 42125
rect 53484 42120 157491 42122
rect 53484 42064 157430 42120
rect 157486 42064 157491 42120
rect 53484 42062 157491 42064
rect 53484 42060 53490 42062
rect 157425 42059 157491 42062
rect 230105 42122 230171 42125
rect 543774 42122 543780 42124
rect 230105 42120 543780 42122
rect 230105 42064 230110 42120
rect 230166 42064 543780 42120
rect 230105 42062 543780 42064
rect 230105 42059 230171 42062
rect 543774 42060 543780 42062
rect 543844 42060 543850 42124
rect 580165 41986 580231 41989
rect 583520 41986 584960 42076
rect 580165 41984 584960 41986
rect 580165 41928 580170 41984
rect 580226 41928 584960 41984
rect 580165 41926 584960 41928
rect 580165 41923 580231 41926
rect 583520 41836 584960 41926
rect 348233 41442 348299 41445
rect 352230 41442 352236 41444
rect 348233 41440 352236 41442
rect 348233 41384 348238 41440
rect 348294 41384 352236 41440
rect 348233 41382 352236 41384
rect 348233 41379 348299 41382
rect 352230 41380 352236 41382
rect 352300 41380 352306 41444
rect 354254 41380 354260 41444
rect 354324 41442 354330 41444
rect 354622 41442 354628 41444
rect 354324 41382 354628 41442
rect 354324 41380 354330 41382
rect 354622 41380 354628 41382
rect 354692 41380 354698 41444
rect 285673 40626 285739 40629
rect 353334 40626 353340 40628
rect 285673 40624 353340 40626
rect 285673 40568 285678 40624
rect 285734 40568 353340 40624
rect 285673 40566 353340 40568
rect 285673 40563 285739 40566
rect 353334 40564 353340 40566
rect 353404 40564 353410 40628
rect 6177 40354 6243 40357
rect 353845 40354 353911 40357
rect 6177 40352 353911 40354
rect 6177 40296 6182 40352
rect 6238 40296 353850 40352
rect 353906 40296 353911 40352
rect 6177 40294 353911 40296
rect 6177 40291 6243 40294
rect 353845 40291 353911 40294
rect 354949 40354 355015 40357
rect 356094 40354 356100 40356
rect 354949 40352 356100 40354
rect 354949 40296 354954 40352
rect 355010 40296 356100 40352
rect 354949 40294 356100 40296
rect 354949 40291 355015 40294
rect 356094 40292 356100 40294
rect 356164 40292 356170 40356
rect 10317 40218 10383 40221
rect 381077 40218 381143 40221
rect 10317 40216 381143 40218
rect 10317 40160 10322 40216
rect 10378 40160 381082 40216
rect 381138 40160 381143 40216
rect 10317 40158 381143 40160
rect 10317 40155 10383 40158
rect 381077 40155 381143 40158
rect 10501 40082 10567 40085
rect 390277 40082 390343 40085
rect 10501 40080 390343 40082
rect 10501 40024 10506 40080
rect 10562 40024 390282 40080
rect 390338 40024 390343 40080
rect 10501 40022 390343 40024
rect 10501 40019 10567 40022
rect 390277 40019 390343 40022
rect 393313 40082 393379 40085
rect 415894 40082 415900 40084
rect 393313 40080 415900 40082
rect 393313 40024 393318 40080
rect 393374 40024 415900 40080
rect 393313 40022 415900 40024
rect 393313 40019 393379 40022
rect 415894 40020 415900 40022
rect 415964 40020 415970 40084
rect 122598 39884 122604 39948
rect 122668 39946 122674 39948
rect 132677 39946 132743 39949
rect 122668 39944 132743 39946
rect 122668 39888 132682 39944
rect 132738 39888 132743 39944
rect 122668 39886 132743 39888
rect 122668 39884 122674 39886
rect 132677 39883 132743 39886
rect 308489 39946 308555 39949
rect 313222 39946 313228 39948
rect 308489 39944 313228 39946
rect 308489 39888 308494 39944
rect 308550 39888 313228 39944
rect 308489 39886 313228 39888
rect 308489 39883 308555 39886
rect 313222 39884 313228 39886
rect 313292 39884 313298 39948
rect 60089 39810 60155 39813
rect 488574 39810 488580 39812
rect 60089 39808 488580 39810
rect 60089 39752 60094 39808
rect 60150 39752 488580 39808
rect 60089 39750 488580 39752
rect 60089 39747 60155 39750
rect 488574 39748 488580 39750
rect 488644 39748 488650 39812
rect 23381 39674 23447 39677
rect 165981 39674 166047 39677
rect 23381 39672 166047 39674
rect 23381 39616 23386 39672
rect 23442 39616 165986 39672
rect 166042 39616 166047 39672
rect 23381 39614 166047 39616
rect 23381 39611 23447 39614
rect 165981 39611 166047 39614
rect 175273 39674 175339 39677
rect 551645 39674 551711 39677
rect 175273 39672 551711 39674
rect 175273 39616 175278 39672
rect 175334 39616 551650 39672
rect 551706 39616 551711 39672
rect 175273 39614 551711 39616
rect 175273 39611 175339 39614
rect 551645 39611 551711 39614
rect 53598 39476 53604 39540
rect 53668 39538 53674 39540
rect 84285 39538 84351 39541
rect 53668 39536 84351 39538
rect 53668 39480 84290 39536
rect 84346 39480 84351 39536
rect 53668 39478 84351 39480
rect 53668 39476 53674 39478
rect 84285 39475 84351 39478
rect 287329 39538 287395 39541
rect 467782 39538 467788 39540
rect 287329 39536 467788 39538
rect 287329 39480 287334 39536
rect 287390 39480 467788 39536
rect 287329 39478 467788 39480
rect 287329 39475 287395 39478
rect 467782 39476 467788 39478
rect 467852 39476 467858 39540
rect 256969 39402 257035 39405
rect 352046 39402 352052 39404
rect 256969 39400 352052 39402
rect -960 39266 480 39356
rect 256969 39344 256974 39400
rect 257030 39344 352052 39400
rect 256969 39342 352052 39344
rect 256969 39339 257035 39342
rect 352046 39340 352052 39342
rect 352116 39340 352122 39404
rect 358670 39340 358676 39404
rect 358740 39402 358746 39404
rect 462957 39402 463023 39405
rect 358740 39400 463023 39402
rect 358740 39344 462962 39400
rect 463018 39344 463023 39400
rect 358740 39342 463023 39344
rect 358740 39340 358746 39342
rect 462957 39339 463023 39342
rect 2773 39266 2839 39269
rect -960 39264 2839 39266
rect -960 39208 2778 39264
rect 2834 39208 2839 39264
rect -960 39206 2839 39208
rect -960 39116 480 39206
rect 2773 39203 2839 39206
rect 317505 39266 317571 39269
rect 365662 39266 365668 39268
rect 317505 39264 365668 39266
rect 317505 39208 317510 39264
rect 317566 39208 365668 39264
rect 317505 39206 365668 39208
rect 317505 39203 317571 39206
rect 365662 39204 365668 39206
rect 365732 39204 365738 39268
rect 350533 39130 350599 39133
rect 353518 39130 353524 39132
rect 350533 39128 353524 39130
rect 350533 39072 350538 39128
rect 350594 39072 353524 39128
rect 350533 39070 353524 39072
rect 350533 39067 350599 39070
rect 353518 39068 353524 39070
rect 353588 39068 353594 39132
rect 367686 39068 367692 39132
rect 367756 39130 367762 39132
rect 423673 39130 423739 39133
rect 367756 39128 423739 39130
rect 367756 39072 423678 39128
rect 423734 39072 423739 39128
rect 367756 39070 423739 39072
rect 367756 39068 367762 39070
rect 423673 39067 423739 39070
rect 3233 38994 3299 38997
rect 471973 38994 472039 38997
rect 3233 38992 472039 38994
rect 3233 38936 3238 38992
rect 3294 38936 471978 38992
rect 472034 38936 472039 38992
rect 3233 38934 472039 38936
rect 3233 38931 3299 38934
rect 471973 38931 472039 38934
rect 362166 38796 362172 38860
rect 362236 38858 362242 38860
rect 432597 38858 432663 38861
rect 362236 38856 432663 38858
rect 362236 38800 432602 38856
rect 432658 38800 432663 38856
rect 362236 38798 432663 38800
rect 362236 38796 362242 38798
rect 432597 38795 432663 38798
rect 364926 38660 364932 38724
rect 364996 38722 365002 38724
rect 378133 38722 378199 38725
rect 364996 38720 378199 38722
rect 364996 38664 378138 38720
rect 378194 38664 378199 38720
rect 364996 38662 378199 38664
rect 364996 38660 365002 38662
rect 378133 38659 378199 38662
rect 580165 37090 580231 37093
rect 583520 37090 584960 37180
rect 580165 37088 584960 37090
rect 580165 37032 580170 37088
rect 580226 37032 584960 37088
rect 580165 37030 584960 37032
rect 580165 37027 580231 37030
rect 583520 36940 584960 37030
rect 354254 35940 354260 36004
rect 354324 36002 354330 36004
rect 354622 36002 354628 36004
rect 354324 35942 354628 36002
rect 354324 35940 354330 35942
rect 354622 35940 354628 35942
rect 354692 35940 354698 36004
rect 354581 35866 354647 35869
rect 354536 35864 354690 35866
rect 354536 35808 354586 35864
rect 354642 35808 354690 35864
rect 354536 35806 354690 35808
rect 354581 35803 354690 35806
rect 354630 35732 354690 35803
rect 354622 35668 354628 35732
rect 354692 35668 354698 35732
rect -960 34370 480 34460
rect 3417 34370 3483 34373
rect -960 34368 3483 34370
rect -960 34312 3422 34368
rect 3478 34312 3483 34368
rect -960 34310 3483 34312
rect -960 34220 480 34310
rect 3417 34307 3483 34310
rect 39062 33764 39068 33828
rect 39132 33826 39138 33828
rect 488533 33826 488599 33829
rect 39132 33824 488599 33826
rect 39132 33768 488538 33824
rect 488594 33768 488599 33824
rect 39132 33766 488599 33768
rect 39132 33764 39138 33766
rect 488533 33763 488599 33766
rect 528553 33826 528619 33829
rect 545062 33826 545068 33828
rect 528553 33824 545068 33826
rect 528553 33768 528558 33824
rect 528614 33768 545068 33824
rect 528553 33766 545068 33768
rect 528553 33763 528619 33766
rect 545062 33764 545068 33766
rect 545132 33764 545138 33828
rect 287697 33554 287763 33557
rect 295926 33554 295932 33556
rect 287697 33552 295932 33554
rect 287697 33496 287702 33552
rect 287758 33496 295932 33552
rect 287697 33494 295932 33496
rect 287697 33491 287763 33494
rect 295926 33492 295932 33494
rect 295996 33492 296002 33556
rect 580073 32194 580139 32197
rect 583520 32194 584960 32284
rect 580073 32192 584960 32194
rect 580073 32136 580078 32192
rect 580134 32136 584960 32192
rect 580073 32134 584960 32136
rect 580073 32131 580139 32134
rect 583520 32044 584960 32134
rect -960 29474 480 29564
rect 3877 29474 3943 29477
rect -960 29472 3943 29474
rect -960 29416 3882 29472
rect 3938 29416 3943 29472
rect -960 29414 3943 29416
rect -960 29324 480 29414
rect 3877 29411 3943 29414
rect 580073 27298 580139 27301
rect 583520 27298 584960 27388
rect 580073 27296 584960 27298
rect 580073 27240 580078 27296
rect 580134 27240 584960 27296
rect 580073 27238 584960 27240
rect 580073 27235 580139 27238
rect 583520 27148 584960 27238
rect 354581 26348 354647 26349
rect 354581 26346 354628 26348
rect 354536 26344 354628 26346
rect 354692 26346 354698 26348
rect 354536 26288 354586 26344
rect 354536 26286 354628 26288
rect 354581 26284 354628 26286
rect 354692 26286 354774 26346
rect 354692 26284 354698 26286
rect 354581 26283 354647 26284
rect 354581 26212 354647 26213
rect 354581 26210 354628 26212
rect 354536 26208 354628 26210
rect 354692 26210 354698 26212
rect 354536 26152 354586 26208
rect 354536 26150 354628 26152
rect 354581 26148 354628 26150
rect 354692 26150 354774 26210
rect 354692 26148 354698 26150
rect 354581 26147 354647 26148
rect -960 24578 480 24668
rect 3233 24578 3299 24581
rect -960 24576 3299 24578
rect -960 24520 3238 24576
rect 3294 24520 3299 24576
rect -960 24518 3299 24520
rect -960 24428 480 24518
rect 3233 24515 3299 24518
rect 580441 22402 580507 22405
rect 583520 22402 584960 22492
rect 580441 22400 584960 22402
rect 580441 22344 580446 22400
rect 580502 22344 584960 22400
rect 580441 22342 584960 22344
rect 580441 22339 580507 22342
rect 583520 22252 584960 22342
rect -960 19682 480 19772
rect 3693 19682 3759 19685
rect -960 19680 3759 19682
rect -960 19624 3698 19680
rect 3754 19624 3759 19680
rect -960 19622 3759 19624
rect -960 19532 480 19622
rect 3693 19619 3759 19622
rect 583520 17506 584960 17596
rect 583342 17446 584960 17506
rect 583342 17370 583402 17446
rect 583520 17370 584960 17446
rect 583342 17356 584960 17370
rect 583342 17310 583586 17356
rect 354581 16690 354647 16693
rect 354806 16690 354812 16692
rect 354536 16688 354812 16690
rect 354536 16632 354586 16688
rect 354642 16632 354812 16688
rect 354536 16630 354812 16632
rect 354581 16627 354647 16630
rect 354806 16628 354812 16630
rect 354876 16628 354882 16692
rect 545614 16628 545620 16692
rect 545684 16690 545690 16692
rect 583526 16690 583586 17310
rect 545684 16630 583586 16690
rect 545684 16628 545690 16630
rect 354581 16556 354647 16557
rect 354581 16554 354628 16556
rect 354536 16552 354628 16554
rect 354692 16554 354698 16556
rect 354536 16496 354586 16552
rect 354536 16494 354628 16496
rect 354581 16492 354628 16494
rect 354692 16494 354774 16554
rect 354692 16492 354698 16494
rect 354581 16491 354647 16492
rect -960 14786 480 14876
rect 3417 14786 3483 14789
rect -960 14784 3483 14786
rect -960 14728 3422 14784
rect 3478 14728 3483 14784
rect -960 14726 3483 14728
rect -960 14636 480 14726
rect 3417 14723 3483 14726
rect 580717 12610 580783 12613
rect 583520 12610 584960 12700
rect 580717 12608 584960 12610
rect 580717 12552 580722 12608
rect 580778 12552 584960 12608
rect 580717 12550 584960 12552
rect 580717 12547 580783 12550
rect 583520 12460 584960 12550
rect 187601 10298 187667 10301
rect 542302 10298 542308 10300
rect 187601 10296 542308 10298
rect 187601 10240 187606 10296
rect 187662 10240 542308 10296
rect 187601 10238 542308 10240
rect 187601 10235 187667 10238
rect 542302 10236 542308 10238
rect 542372 10236 542378 10300
rect -960 9890 480 9980
rect 2957 9890 3023 9893
rect -960 9888 3023 9890
rect -960 9832 2962 9888
rect 3018 9832 3023 9888
rect -960 9830 3023 9832
rect -960 9740 480 9830
rect 2957 9827 3023 9830
rect 207606 8876 207612 8940
rect 207676 8938 207682 8940
rect 213821 8938 213887 8941
rect 207676 8936 213887 8938
rect 207676 8880 213826 8936
rect 213882 8880 213887 8936
rect 207676 8878 213887 8880
rect 207676 8876 207682 8878
rect 213821 8875 213887 8878
rect 580165 7714 580231 7717
rect 583520 7714 584960 7804
rect 580165 7712 584960 7714
rect 580165 7656 580170 7712
rect 580226 7656 584960 7712
rect 580165 7654 584960 7656
rect 580165 7651 580231 7654
rect 583520 7564 584960 7654
rect 354622 7108 354628 7172
rect 354692 7108 354698 7172
rect 354630 7037 354690 7108
rect 354581 7034 354690 7037
rect 354536 7032 354690 7034
rect 354536 6976 354586 7032
rect 354642 6976 354690 7032
rect 354536 6974 354690 6976
rect 354581 6971 354647 6974
rect 309501 6490 309567 6493
rect 443494 6490 443500 6492
rect 309501 6488 443500 6490
rect 309501 6432 309506 6488
rect 309562 6432 443500 6488
rect 309501 6430 443500 6432
rect 309501 6427 309567 6430
rect 443494 6428 443500 6430
rect 443564 6428 443570 6492
rect 246205 6354 246271 6357
rect 541014 6354 541020 6356
rect 246205 6352 541020 6354
rect 246205 6296 246210 6352
rect 246266 6296 541020 6352
rect 246205 6294 541020 6296
rect 246205 6291 246271 6294
rect 541014 6292 541020 6294
rect 541084 6292 541090 6356
rect 83181 6218 83247 6221
rect 541198 6218 541204 6220
rect 83181 6216 541204 6218
rect 83181 6160 83186 6216
rect 83242 6160 541204 6216
rect 83181 6158 541204 6160
rect 83181 6155 83247 6158
rect 541198 6156 541204 6158
rect 541268 6156 541274 6220
rect 302877 5538 302943 5541
rect 394734 5538 394740 5540
rect 302877 5536 394740 5538
rect 302877 5480 302882 5536
rect 302938 5480 394740 5536
rect 302877 5478 394740 5480
rect 302877 5475 302943 5478
rect 394734 5476 394740 5478
rect 394804 5476 394810 5540
rect 99741 5402 99807 5405
rect 354438 5402 354444 5404
rect 99741 5400 354444 5402
rect 99741 5344 99746 5400
rect 99802 5344 354444 5400
rect 99741 5342 354444 5344
rect 99741 5339 99807 5342
rect 354438 5340 354444 5342
rect 354508 5340 354514 5404
rect 239581 5266 239647 5269
rect 524454 5266 524460 5268
rect 239581 5264 524460 5266
rect 239581 5208 239586 5264
rect 239642 5208 524460 5264
rect 239581 5206 524460 5208
rect 239581 5203 239647 5206
rect 524454 5204 524460 5206
rect 524524 5204 524530 5268
rect 209589 5130 209655 5133
rect 545246 5130 545252 5132
rect 209589 5128 545252 5130
rect -960 4994 480 5084
rect 209589 5072 209594 5128
rect 209650 5072 545252 5128
rect 209589 5070 545252 5072
rect 209589 5067 209655 5070
rect 545246 5068 545252 5070
rect 545316 5068 545322 5132
rect 2773 4994 2839 4997
rect -960 4992 2839 4994
rect -960 4936 2778 4992
rect 2834 4936 2839 4992
rect -960 4934 2839 4936
rect -960 4844 480 4934
rect 2773 4931 2839 4934
rect 39798 4932 39804 4996
rect 39868 4994 39874 4996
rect 419349 4994 419415 4997
rect 39868 4992 419415 4994
rect 39868 4936 419354 4992
rect 419410 4936 419415 4992
rect 39868 4934 419415 4936
rect 39868 4932 39874 4934
rect 419349 4931 419415 4934
rect 476021 4994 476087 4997
rect 512126 4994 512132 4996
rect 476021 4992 512132 4994
rect 476021 4936 476026 4992
rect 476082 4936 512132 4992
rect 476021 4934 512132 4936
rect 476021 4931 476087 4934
rect 512126 4932 512132 4934
rect 512196 4932 512202 4996
rect 96429 4858 96495 4861
rect 543958 4858 543964 4860
rect 96429 4856 543964 4858
rect 96429 4800 96434 4856
rect 96490 4800 543964 4856
rect 96429 4798 543964 4800
rect 96429 4795 96495 4798
rect 543958 4796 543964 4798
rect 544028 4796 544034 4860
rect 42374 3980 42380 4044
rect 42444 4042 42450 4044
rect 202965 4042 203031 4045
rect 42444 4040 203031 4042
rect 42444 3984 202970 4040
rect 203026 3984 203031 4040
rect 42444 3982 203031 3984
rect 42444 3980 42450 3982
rect 202965 3979 203031 3982
rect 249517 4042 249583 4045
rect 466494 4042 466500 4044
rect 249517 4040 466500 4042
rect 249517 3984 249522 4040
rect 249578 3984 466500 4040
rect 249517 3982 466500 3984
rect 249517 3979 249583 3982
rect 466494 3980 466500 3982
rect 466564 3980 466570 4044
rect 55070 3844 55076 3908
rect 55140 3906 55146 3908
rect 339493 3906 339559 3909
rect 55140 3904 339559 3906
rect 55140 3848 339498 3904
rect 339554 3848 339559 3904
rect 55140 3846 339559 3848
rect 55140 3844 55146 3846
rect 339493 3843 339559 3846
rect 358854 3844 358860 3908
rect 358924 3906 358930 3908
rect 359365 3906 359431 3909
rect 358924 3904 359431 3906
rect 358924 3848 359370 3904
rect 359426 3848 359431 3904
rect 358924 3846 359431 3848
rect 358924 3844 358930 3846
rect 359365 3843 359431 3846
rect 368974 3844 368980 3908
rect 369044 3906 369050 3908
rect 519261 3906 519327 3909
rect 369044 3904 519327 3906
rect 369044 3848 519266 3904
rect 519322 3848 519327 3904
rect 369044 3846 519327 3848
rect 369044 3844 369050 3846
rect 519261 3843 519327 3846
rect 116485 3770 116551 3773
rect 451038 3770 451044 3772
rect 116485 3768 451044 3770
rect 116485 3712 116490 3768
rect 116546 3712 451044 3768
rect 116485 3710 451044 3712
rect 116485 3707 116551 3710
rect 451038 3708 451044 3710
rect 451108 3708 451114 3772
rect 73245 3634 73311 3637
rect 460974 3634 460980 3636
rect 73245 3632 460980 3634
rect 73245 3576 73250 3632
rect 73306 3576 460980 3632
rect 73245 3574 460980 3576
rect 73245 3571 73311 3574
rect 460974 3572 460980 3574
rect 461044 3572 461050 3636
rect 515254 3572 515260 3636
rect 515324 3634 515330 3636
rect 515949 3634 516015 3637
rect 515324 3632 516015 3634
rect 515324 3576 515954 3632
rect 516010 3576 516015 3632
rect 515324 3574 516015 3576
rect 515324 3572 515330 3574
rect 515949 3571 516015 3574
rect 42558 3436 42564 3500
rect 42628 3498 42634 3500
rect 56501 3498 56567 3501
rect 42628 3496 56567 3498
rect 42628 3440 56506 3496
rect 56562 3440 56567 3496
rect 42628 3438 56567 3440
rect 42628 3436 42634 3438
rect 56501 3435 56567 3438
rect 106365 3498 106431 3501
rect 543038 3498 543044 3500
rect 106365 3496 543044 3498
rect 106365 3440 106370 3496
rect 106426 3440 543044 3496
rect 106365 3438 543044 3440
rect 106365 3435 106431 3438
rect 543038 3436 543044 3438
rect 543108 3436 543114 3500
rect 39246 3300 39252 3364
rect 39316 3362 39322 3364
rect 479333 3362 479399 3365
rect 39316 3360 479399 3362
rect 39316 3304 479338 3360
rect 479394 3304 479399 3360
rect 39316 3302 479399 3304
rect 39316 3300 39322 3302
rect 479333 3299 479399 3302
rect 354254 3164 354260 3228
rect 354324 3226 354330 3228
rect 439405 3226 439471 3229
rect 354324 3224 439471 3226
rect 354324 3168 439410 3224
rect 439466 3168 439471 3224
rect 354324 3166 439471 3168
rect 354324 3164 354330 3166
rect 439405 3163 439471 3166
rect 356646 3028 356652 3092
rect 356716 3090 356722 3092
rect 362677 3090 362743 3093
rect 356716 3088 362743 3090
rect 356716 3032 362682 3088
rect 362738 3032 362743 3088
rect 356716 3030 362743 3032
rect 356716 3028 356722 3030
rect 362677 3027 362743 3030
rect 363454 3028 363460 3092
rect 363524 3090 363530 3092
rect 412725 3090 412791 3093
rect 363524 3088 412791 3090
rect 363524 3032 412730 3088
rect 412786 3032 412791 3088
rect 363524 3030 412791 3032
rect 363524 3028 363530 3030
rect 412725 3027 412791 3030
rect 425094 3028 425100 3092
rect 425164 3090 425170 3092
rect 425973 3090 426039 3093
rect 425164 3088 426039 3090
rect 425164 3032 425978 3088
rect 426034 3032 426039 3088
rect 425164 3030 426039 3032
rect 425164 3028 425170 3030
rect 425973 3027 426039 3030
rect 432597 3090 432663 3093
rect 440182 3090 440188 3092
rect 432597 3088 440188 3090
rect 432597 3032 432602 3088
rect 432658 3032 440188 3088
rect 432597 3030 440188 3032
rect 432597 3027 432663 3030
rect 440182 3028 440188 3030
rect 440252 3028 440258 3092
rect 459277 3090 459343 3093
rect 441570 3088 459343 3090
rect 441570 3032 459282 3088
rect 459338 3032 459343 3088
rect 441570 3030 459343 3032
rect 360694 2892 360700 2956
rect 360764 2954 360770 2956
rect 392669 2954 392735 2957
rect 402789 2956 402855 2957
rect 402789 2954 402836 2956
rect 360764 2952 392735 2954
rect 360764 2896 392674 2952
rect 392730 2896 392735 2952
rect 360764 2894 392735 2896
rect 402744 2952 402836 2954
rect 402744 2896 402794 2952
rect 402744 2894 402836 2896
rect 360764 2892 360770 2894
rect 392669 2891 392735 2894
rect 402789 2892 402836 2894
rect 402900 2892 402906 2956
rect 436686 2892 436692 2956
rect 436756 2954 436762 2956
rect 441570 2954 441630 3030
rect 459277 3027 459343 3030
rect 436756 2894 441630 2954
rect 436756 2892 436762 2894
rect 402789 2891 402855 2892
rect 580165 2818 580231 2821
rect 583520 2818 584960 2908
rect 580165 2816 584960 2818
rect 580165 2760 580170 2816
rect 580226 2760 584960 2816
rect 580165 2758 584960 2760
rect 580165 2755 580231 2758
rect 583520 2668 584960 2758
<< via3 >>
rect 541940 700980 542004 701044
rect 39620 700844 39684 700908
rect 405596 700844 405660 700908
rect 39068 700708 39132 700772
rect 542860 700572 542924 700636
rect 542492 700436 542556 700500
rect 40540 700300 40604 700364
rect 370452 700164 370516 700228
rect 415900 700164 415964 700228
rect 362172 700028 362236 700092
rect 59860 699892 59924 699956
rect 39988 699756 40052 699820
rect 364932 699892 364996 699956
rect 66300 699816 66364 699820
rect 66300 699760 66314 699816
rect 66314 699760 66364 699816
rect 66300 699756 66364 699760
rect 333836 699756 333900 699820
rect 367692 699892 367756 699956
rect 365668 699756 365732 699820
rect 467788 699756 467852 699820
rect 488580 699756 488644 699820
rect 543780 699756 543844 699820
rect 353340 668476 353404 668540
rect 55996 666436 56060 666500
rect 351868 666436 351932 666500
rect 368980 664668 369044 664732
rect 363460 664532 363524 664596
rect 42748 664396 42812 664460
rect 436692 664396 436756 664460
rect 55076 664260 55140 664324
rect 360700 664260 360764 664324
rect 402836 664260 402900 664324
rect 545068 664124 545132 664188
rect 42380 663988 42444 664052
rect 310468 663852 310532 663916
rect 443500 663852 443564 663916
rect 541020 663852 541084 663916
rect 354812 663716 354876 663780
rect 59860 662688 59924 662692
rect 59860 662632 59910 662688
rect 59910 662632 59924 662688
rect 59860 662628 59924 662632
rect 355364 662356 355428 662420
rect 285812 662084 285876 662148
rect 297956 662084 298020 662148
rect 301452 662144 301516 662148
rect 301452 662088 301466 662144
rect 301466 662088 301516 662144
rect 301452 662084 301516 662088
rect 53236 661948 53300 662012
rect 98684 661948 98748 662012
rect 172468 661948 172532 662012
rect 356100 662220 356164 662284
rect 354076 662144 354140 662148
rect 354076 662088 354090 662144
rect 354090 662088 354140 662144
rect 354076 662084 354140 662088
rect 358676 662084 358740 662148
rect 354444 661948 354508 662012
rect 53420 661812 53484 661876
rect 179460 661872 179524 661876
rect 179460 661816 179510 661872
rect 179510 661816 179524 661872
rect 179460 661812 179524 661816
rect 358860 661948 358924 662012
rect 356652 661812 356716 661876
rect 366036 661812 366100 661876
rect 394740 661872 394804 661876
rect 394740 661816 394790 661872
rect 394790 661816 394804 661872
rect 394740 661812 394804 661816
rect 440188 661872 440252 661876
rect 440188 661816 440238 661872
rect 440238 661816 440252 661872
rect 440188 661812 440252 661816
rect 451044 661812 451108 661876
rect 460980 661812 461044 661876
rect 466500 661812 466564 661876
rect 38884 661676 38948 661740
rect 512132 661676 512196 661740
rect 515260 661736 515324 661740
rect 515260 661680 515274 661736
rect 515274 661680 515324 661736
rect 515260 661676 515324 661680
rect 524460 661676 524524 661740
rect 121500 661540 121564 661604
rect 108988 661404 109052 661468
rect 49740 661268 49804 661332
rect 541756 661268 541820 661332
rect 366036 661132 366100 661196
rect 98684 660996 98748 661060
rect 545620 660996 545684 661060
rect 53604 660860 53668 660924
rect 66300 660860 66364 660924
rect 333836 660860 333900 660924
rect 352052 660860 352116 660924
rect 544332 660860 544396 660924
rect 108988 660724 109052 660788
rect 310468 660724 310532 660788
rect 352236 660724 352300 660788
rect 121500 660588 121564 660652
rect 301452 660588 301516 660652
rect 353524 660588 353588 660652
rect 46244 660452 46308 660516
rect 54708 660452 54772 660516
rect 172468 660452 172532 660516
rect 285812 660452 285876 660516
rect 352420 660452 352484 660516
rect 543596 660452 543660 660516
rect 49740 660316 49804 660380
rect 54892 660316 54956 660380
rect 179460 660316 179524 660380
rect 297956 660316 298020 660380
rect 425100 660316 425164 660380
rect 544516 660316 544580 660380
rect 542124 660180 542188 660244
rect 542308 660180 542372 660244
rect 46244 659908 46308 659972
rect 39252 657384 39316 657388
rect 39252 657328 39302 657384
rect 39302 657328 39316 657384
rect 39252 657324 39316 657328
rect 542124 653380 542188 653444
rect 39804 623732 39868 623796
rect 39436 610404 39500 610468
rect 39252 606188 39316 606252
rect 542308 592860 542372 592924
rect 542308 587692 542372 587756
rect 545252 583204 545316 583268
rect 40540 582388 40604 582452
rect 543964 542948 544028 543012
rect 39252 516292 39316 516356
rect 542124 482156 542188 482220
rect 541940 471880 542004 471884
rect 541940 471824 541990 471880
rect 541990 471824 542004 471880
rect 541940 471820 542004 471824
rect 544148 471412 544212 471476
rect 541756 468284 541820 468348
rect 541756 468012 541820 468076
rect 541940 466304 542004 466308
rect 541940 466248 541990 466304
rect 541990 466248 542004 466304
rect 541940 466244 542004 466248
rect 541940 445708 542004 445772
rect 541756 444348 541820 444412
rect 541756 442444 541820 442508
rect 541756 439044 541820 439108
rect 541756 438908 541820 438972
rect 541756 438092 541820 438156
rect 40172 404500 40236 404564
rect 39068 382332 39132 382396
rect 543044 369140 543108 369204
rect 39068 364380 39132 364444
rect 38884 359756 38948 359820
rect 38884 337316 38948 337380
rect 542676 296652 542740 296716
rect 541756 291076 541820 291140
rect 542492 284140 542556 284204
rect 544516 261020 544580 261084
rect 544332 234092 544396 234156
rect 543596 191660 543660 191724
rect 541756 150452 541820 150516
rect 542860 139436 542924 139500
rect 544332 135492 544396 135556
rect 39620 117948 39684 118012
rect 39988 55388 40052 55452
rect 541940 49540 542004 49604
rect 544332 49540 544396 49604
rect 40172 44644 40236 44708
rect 542676 44508 542740 44572
rect 541756 44372 541820 44436
rect 541572 44236 541636 44300
rect 38884 44100 38948 44164
rect 541940 43964 542004 44028
rect 55996 43828 56060 43892
rect 122604 43828 122668 43892
rect 283972 43828 284036 43892
rect 354812 43828 354876 43892
rect 53236 43692 53300 43756
rect 207612 43692 207676 43756
rect 223988 43692 224052 43756
rect 351868 43692 351932 43756
rect 39436 43556 39500 43620
rect 544148 43420 544212 43484
rect 295932 43284 295996 43348
rect 355180 43284 355244 43348
rect 313228 43148 313292 43212
rect 352420 43148 352484 43212
rect 54892 42332 54956 42396
rect 223988 42392 224052 42396
rect 223988 42336 224002 42392
rect 224002 42336 224052 42392
rect 223988 42332 224052 42336
rect 283972 42392 284036 42396
rect 283972 42336 284022 42392
rect 284022 42336 284036 42392
rect 283972 42332 284036 42336
rect 370452 42332 370516 42396
rect 405596 42392 405660 42396
rect 405596 42336 405610 42392
rect 405610 42336 405660 42392
rect 405596 42332 405660 42336
rect 54708 42196 54772 42260
rect 53420 42060 53484 42124
rect 543780 42060 543844 42124
rect 352236 41380 352300 41444
rect 354260 41380 354324 41444
rect 354628 41380 354692 41444
rect 353340 40564 353404 40628
rect 356100 40292 356164 40356
rect 415900 40020 415964 40084
rect 122604 39884 122668 39948
rect 313228 39884 313292 39948
rect 488580 39748 488644 39812
rect 53604 39476 53668 39540
rect 467788 39476 467852 39540
rect 352052 39340 352116 39404
rect 358676 39340 358740 39404
rect 365668 39204 365732 39268
rect 353524 39068 353588 39132
rect 367692 39068 367756 39132
rect 362172 38796 362236 38860
rect 364932 38660 364996 38724
rect 354260 35940 354324 36004
rect 354628 35940 354692 36004
rect 354628 35668 354692 35732
rect 39068 33764 39132 33828
rect 545068 33764 545132 33828
rect 295932 33492 295996 33556
rect 354628 26344 354692 26348
rect 354628 26288 354642 26344
rect 354642 26288 354692 26344
rect 354628 26284 354692 26288
rect 354628 26208 354692 26212
rect 354628 26152 354642 26208
rect 354642 26152 354692 26208
rect 354628 26148 354692 26152
rect 354812 16628 354876 16692
rect 545620 16628 545684 16692
rect 354628 16552 354692 16556
rect 354628 16496 354642 16552
rect 354642 16496 354692 16552
rect 354628 16492 354692 16496
rect 542308 10236 542372 10300
rect 207612 8876 207676 8940
rect 354628 7108 354692 7172
rect 443500 6428 443564 6492
rect 541020 6292 541084 6356
rect 541204 6156 541268 6220
rect 394740 5476 394804 5540
rect 354444 5340 354508 5404
rect 524460 5204 524524 5268
rect 545252 5068 545316 5132
rect 39804 4932 39868 4996
rect 512132 4932 512196 4996
rect 543964 4796 544028 4860
rect 42380 3980 42444 4044
rect 466500 3980 466564 4044
rect 55076 3844 55140 3908
rect 358860 3844 358924 3908
rect 368980 3844 369044 3908
rect 451044 3708 451108 3772
rect 460980 3572 461044 3636
rect 515260 3572 515324 3636
rect 42564 3436 42628 3500
rect 543044 3436 543108 3500
rect 39252 3300 39316 3364
rect 354260 3164 354324 3228
rect 356652 3028 356716 3092
rect 363460 3028 363524 3092
rect 425100 3028 425164 3092
rect 440188 3028 440252 3092
rect 360700 2892 360764 2956
rect 402836 2952 402900 2956
rect 402836 2896 402850 2952
rect 402850 2896 402900 2952
rect 402836 2892 402900 2896
rect 436692 2892 436756 2956
<< metal4 >>
rect 541939 701044 542005 701045
rect 541939 700980 541940 701044
rect 542004 700980 542005 701044
rect 541939 700979 542005 700980
rect 39619 700908 39685 700909
rect 39619 700844 39620 700908
rect 39684 700844 39685 700908
rect 39619 700843 39685 700844
rect 405595 700908 405661 700909
rect 405595 700844 405596 700908
rect 405660 700844 405661 700908
rect 405595 700843 405661 700844
rect 39067 700772 39133 700773
rect 39067 700708 39068 700772
rect 39132 700708 39133 700772
rect 39067 700707 39133 700708
rect 38883 661740 38949 661741
rect 38883 661676 38884 661740
rect 38948 661676 38949 661740
rect 38883 661675 38949 661676
rect 38886 359821 38946 661675
rect 39070 382397 39130 700707
rect 39251 657388 39317 657389
rect 39251 657324 39252 657388
rect 39316 657324 39317 657388
rect 39251 657323 39317 657324
rect 39254 606253 39314 657323
rect 39435 610468 39501 610469
rect 39435 610404 39436 610468
rect 39500 610404 39501 610468
rect 39435 610403 39501 610404
rect 39251 606252 39317 606253
rect 39251 606188 39252 606252
rect 39316 606188 39317 606252
rect 39251 606187 39317 606188
rect 39251 516356 39317 516357
rect 39251 516292 39252 516356
rect 39316 516292 39317 516356
rect 39251 516291 39317 516292
rect 39067 382396 39133 382397
rect 39067 382332 39068 382396
rect 39132 382332 39133 382396
rect 39067 382331 39133 382332
rect 39067 364444 39133 364445
rect 39067 364380 39068 364444
rect 39132 364380 39133 364444
rect 39067 364379 39133 364380
rect 38883 359820 38949 359821
rect 38883 359756 38884 359820
rect 38948 359756 38949 359820
rect 38883 359755 38949 359756
rect 38883 337380 38949 337381
rect 38883 337316 38884 337380
rect 38948 337316 38949 337380
rect 38883 337315 38949 337316
rect 38886 44165 38946 337315
rect 38883 44164 38949 44165
rect 38883 44100 38884 44164
rect 38948 44100 38949 44164
rect 38883 44099 38949 44100
rect 39070 33829 39130 364379
rect 39067 33828 39133 33829
rect 39067 33764 39068 33828
rect 39132 33764 39133 33828
rect 39067 33763 39133 33764
rect 39254 3365 39314 516291
rect 39438 43621 39498 610403
rect 39622 118013 39682 700843
rect 40539 700364 40605 700365
rect 40539 700300 40540 700364
rect 40604 700300 40605 700364
rect 40539 700299 40605 700300
rect 39987 699820 40053 699821
rect 39987 699756 39988 699820
rect 40052 699756 40053 699820
rect 39987 699755 40053 699756
rect 39803 623796 39869 623797
rect 39803 623732 39804 623796
rect 39868 623732 39869 623796
rect 39803 623731 39869 623732
rect 39619 118012 39685 118013
rect 39619 117948 39620 118012
rect 39684 117948 39685 118012
rect 39619 117947 39685 117948
rect 39435 43620 39501 43621
rect 39435 43556 39436 43620
rect 39500 43556 39501 43620
rect 39435 43555 39501 43556
rect 39806 4997 39866 623731
rect 39990 55453 40050 699755
rect 40542 582453 40602 700299
rect 370451 700228 370517 700229
rect 370451 700164 370452 700228
rect 370516 700164 370517 700228
rect 370451 700163 370517 700164
rect 362171 700092 362237 700093
rect 362171 700028 362172 700092
rect 362236 700028 362237 700092
rect 362171 700027 362237 700028
rect 59859 699956 59925 699957
rect 59859 699892 59860 699956
rect 59924 699892 59925 699956
rect 59859 699891 59925 699892
rect 55995 666500 56061 666501
rect 55995 666436 55996 666500
rect 56060 666436 56061 666500
rect 55995 666435 56061 666436
rect 42747 664460 42813 664461
rect 42747 664396 42748 664460
rect 42812 664396 42813 664460
rect 42747 664395 42813 664396
rect 42379 664052 42445 664053
rect 42379 663988 42380 664052
rect 42444 663988 42445 664052
rect 42379 663987 42445 663988
rect 40539 582452 40605 582453
rect 40539 582388 40540 582452
rect 40604 582388 40605 582452
rect 40539 582387 40605 582388
rect 40171 404564 40237 404565
rect 40171 404500 40172 404564
rect 40236 404500 40237 404564
rect 40171 404499 40237 404500
rect 39987 55452 40053 55453
rect 39987 55388 39988 55452
rect 40052 55388 40053 55452
rect 39987 55387 40053 55388
rect 40174 44709 40234 404499
rect 40171 44708 40237 44709
rect 40171 44644 40172 44708
rect 40236 44644 40237 44708
rect 40171 44643 40237 44644
rect 39803 4996 39869 4997
rect 39803 4932 39804 4996
rect 39868 4932 39869 4996
rect 39803 4931 39869 4932
rect 42382 4045 42442 663987
rect 42750 644490 42810 664395
rect 55075 664324 55141 664325
rect 55075 664260 55076 664324
rect 55140 664260 55141 664324
rect 55075 664259 55141 664260
rect 53235 662012 53301 662013
rect 53235 661948 53236 662012
rect 53300 661948 53301 662012
rect 53235 661947 53301 661948
rect 49739 661332 49805 661333
rect 49739 661268 49740 661332
rect 49804 661268 49805 661332
rect 49739 661267 49805 661268
rect 46243 660516 46309 660517
rect 46243 660452 46244 660516
rect 46308 660452 46309 660516
rect 46243 660451 46309 660452
rect 46246 659973 46306 660451
rect 49742 660381 49802 661267
rect 49739 660380 49805 660381
rect 49739 660316 49740 660380
rect 49804 660316 49805 660380
rect 49739 660315 49805 660316
rect 46243 659972 46309 659973
rect 46243 659908 46244 659972
rect 46308 659908 46309 659972
rect 46243 659907 46309 659908
rect 42566 644430 42810 644490
rect 42379 4044 42445 4045
rect 42379 3980 42380 4044
rect 42444 3980 42445 4044
rect 42379 3979 42445 3980
rect 42566 3501 42626 644430
rect 53238 43757 53298 661947
rect 53419 661876 53485 661877
rect 53419 661812 53420 661876
rect 53484 661812 53485 661876
rect 53419 661811 53485 661812
rect 53235 43756 53301 43757
rect 53235 43692 53236 43756
rect 53300 43692 53301 43756
rect 53235 43691 53301 43692
rect 53422 42125 53482 661811
rect 53603 660924 53669 660925
rect 53603 660860 53604 660924
rect 53668 660860 53669 660924
rect 53603 660859 53669 660860
rect 53419 42124 53485 42125
rect 53419 42060 53420 42124
rect 53484 42060 53485 42124
rect 53419 42059 53485 42060
rect 53606 39541 53666 660859
rect 54707 660516 54773 660517
rect 54707 660452 54708 660516
rect 54772 660452 54773 660516
rect 54707 660451 54773 660452
rect 54710 42261 54770 660451
rect 54891 660380 54957 660381
rect 54891 660316 54892 660380
rect 54956 660316 54957 660380
rect 54891 660315 54957 660316
rect 54894 42397 54954 660315
rect 54891 42396 54957 42397
rect 54891 42332 54892 42396
rect 54956 42332 54957 42396
rect 54891 42331 54957 42332
rect 54707 42260 54773 42261
rect 54707 42196 54708 42260
rect 54772 42196 54773 42260
rect 54707 42195 54773 42196
rect 53603 39540 53669 39541
rect 53603 39476 53604 39540
rect 53668 39476 53669 39540
rect 53603 39475 53669 39476
rect 55078 3909 55138 664259
rect 55998 43893 56058 666435
rect 59862 662693 59922 699891
rect 66299 699820 66365 699821
rect 66299 699756 66300 699820
rect 66364 699756 66365 699820
rect 66299 699755 66365 699756
rect 333835 699820 333901 699821
rect 333835 699756 333836 699820
rect 333900 699756 333901 699820
rect 333835 699755 333901 699756
rect 59859 662692 59925 662693
rect 59859 662628 59860 662692
rect 59924 662628 59925 662692
rect 59859 662627 59925 662628
rect 66302 660925 66362 699755
rect 310467 663916 310533 663917
rect 310467 663852 310468 663916
rect 310532 663852 310533 663916
rect 310467 663851 310533 663852
rect 285811 662148 285877 662149
rect 285811 662084 285812 662148
rect 285876 662084 285877 662148
rect 285811 662083 285877 662084
rect 297955 662148 298021 662149
rect 297955 662084 297956 662148
rect 298020 662084 298021 662148
rect 297955 662083 298021 662084
rect 301451 662148 301517 662149
rect 301451 662084 301452 662148
rect 301516 662084 301517 662148
rect 301451 662083 301517 662084
rect 98683 662012 98749 662013
rect 98683 661948 98684 662012
rect 98748 661948 98749 662012
rect 98683 661947 98749 661948
rect 172467 662012 172533 662013
rect 172467 661948 172468 662012
rect 172532 661948 172533 662012
rect 172467 661947 172533 661948
rect 98686 661061 98746 661947
rect 121499 661604 121565 661605
rect 121499 661540 121500 661604
rect 121564 661540 121565 661604
rect 121499 661539 121565 661540
rect 108987 661468 109053 661469
rect 108987 661404 108988 661468
rect 109052 661404 109053 661468
rect 108987 661403 109053 661404
rect 98683 661060 98749 661061
rect 98683 660996 98684 661060
rect 98748 660996 98749 661060
rect 98683 660995 98749 660996
rect 66299 660924 66365 660925
rect 66299 660860 66300 660924
rect 66364 660860 66365 660924
rect 66299 660859 66365 660860
rect 108990 660789 109050 661403
rect 108987 660788 109053 660789
rect 108987 660724 108988 660788
rect 109052 660724 109053 660788
rect 108987 660723 109053 660724
rect 121502 660653 121562 661539
rect 121499 660652 121565 660653
rect 121499 660588 121500 660652
rect 121564 660588 121565 660652
rect 121499 660587 121565 660588
rect 172470 660517 172530 661947
rect 179459 661876 179525 661877
rect 179459 661812 179460 661876
rect 179524 661812 179525 661876
rect 179459 661811 179525 661812
rect 172467 660516 172533 660517
rect 172467 660452 172468 660516
rect 172532 660452 172533 660516
rect 172467 660451 172533 660452
rect 179462 660381 179522 661811
rect 285814 660517 285874 662083
rect 285811 660516 285877 660517
rect 285811 660452 285812 660516
rect 285876 660452 285877 660516
rect 285811 660451 285877 660452
rect 297958 660381 298018 662083
rect 301454 660653 301514 662083
rect 310470 660789 310530 663851
rect 333838 660925 333898 699755
rect 353339 668540 353405 668541
rect 353339 668476 353340 668540
rect 353404 668476 353405 668540
rect 353339 668475 353405 668476
rect 351867 666500 351933 666501
rect 351867 666436 351868 666500
rect 351932 666436 351933 666500
rect 351867 666435 351933 666436
rect 333835 660924 333901 660925
rect 333835 660860 333836 660924
rect 333900 660860 333901 660924
rect 333835 660859 333901 660860
rect 310467 660788 310533 660789
rect 310467 660724 310468 660788
rect 310532 660724 310533 660788
rect 310467 660723 310533 660724
rect 301451 660652 301517 660653
rect 301451 660588 301452 660652
rect 301516 660588 301517 660652
rect 301451 660587 301517 660588
rect 179459 660380 179525 660381
rect 179459 660316 179460 660380
rect 179524 660316 179525 660380
rect 179459 660315 179525 660316
rect 297955 660380 298021 660381
rect 297955 660316 297956 660380
rect 298020 660316 298021 660380
rect 297955 660315 298021 660316
rect 55995 43892 56061 43893
rect 55995 43828 55996 43892
rect 56060 43828 56061 43892
rect 55995 43827 56061 43828
rect 122603 43892 122669 43893
rect 122603 43828 122604 43892
rect 122668 43828 122669 43892
rect 122603 43827 122669 43828
rect 283971 43892 284037 43893
rect 283971 43828 283972 43892
rect 284036 43828 284037 43892
rect 283971 43827 284037 43828
rect 122606 39949 122666 43827
rect 207611 43756 207677 43757
rect 207611 43692 207612 43756
rect 207676 43692 207677 43756
rect 207611 43691 207677 43692
rect 223987 43756 224053 43757
rect 223987 43692 223988 43756
rect 224052 43692 224053 43756
rect 223987 43691 224053 43692
rect 122603 39948 122669 39949
rect 122603 39884 122604 39948
rect 122668 39884 122669 39948
rect 122603 39883 122669 39884
rect 207614 8941 207674 43691
rect 223990 42397 224050 43691
rect 283974 42397 284034 43827
rect 351870 43757 351930 666435
rect 352051 660924 352117 660925
rect 352051 660860 352052 660924
rect 352116 660860 352117 660924
rect 352051 660859 352117 660860
rect 351867 43756 351933 43757
rect 351867 43692 351868 43756
rect 351932 43692 351933 43756
rect 351867 43691 351933 43692
rect 295931 43348 295997 43349
rect 295931 43284 295932 43348
rect 295996 43284 295997 43348
rect 295931 43283 295997 43284
rect 223987 42396 224053 42397
rect 223987 42332 223988 42396
rect 224052 42332 224053 42396
rect 223987 42331 224053 42332
rect 283971 42396 284037 42397
rect 283971 42332 283972 42396
rect 284036 42332 284037 42396
rect 283971 42331 284037 42332
rect 295934 33557 295994 43283
rect 313227 43212 313293 43213
rect 313227 43148 313228 43212
rect 313292 43148 313293 43212
rect 313227 43147 313293 43148
rect 313230 39949 313290 43147
rect 313227 39948 313293 39949
rect 313227 39884 313228 39948
rect 313292 39884 313293 39948
rect 313227 39883 313293 39884
rect 352054 39405 352114 660859
rect 352235 660788 352301 660789
rect 352235 660724 352236 660788
rect 352300 660724 352301 660788
rect 352235 660723 352301 660724
rect 352238 41445 352298 660723
rect 352419 660516 352485 660517
rect 352419 660452 352420 660516
rect 352484 660452 352485 660516
rect 352419 660451 352485 660452
rect 352422 43213 352482 660451
rect 352419 43212 352485 43213
rect 352419 43148 352420 43212
rect 352484 43148 352485 43212
rect 352419 43147 352485 43148
rect 352235 41444 352301 41445
rect 352235 41380 352236 41444
rect 352300 41380 352301 41444
rect 352235 41379 352301 41380
rect 353342 40629 353402 668475
rect 360699 664324 360765 664325
rect 360699 664260 360700 664324
rect 360764 664260 360765 664324
rect 360699 664259 360765 664260
rect 354811 663780 354877 663781
rect 354811 663716 354812 663780
rect 354876 663716 354877 663780
rect 354811 663715 354877 663716
rect 354075 662148 354141 662149
rect 354075 662084 354076 662148
rect 354140 662084 354141 662148
rect 354075 662083 354141 662084
rect 353523 660652 353589 660653
rect 353523 660588 353524 660652
rect 353588 660588 353589 660652
rect 353523 660587 353589 660588
rect 353339 40628 353405 40629
rect 353339 40564 353340 40628
rect 353404 40564 353405 40628
rect 353339 40563 353405 40564
rect 352051 39404 352117 39405
rect 352051 39340 352052 39404
rect 352116 39340 352117 39404
rect 352051 39339 352117 39340
rect 353526 39133 353586 660587
rect 354078 654150 354138 662083
rect 354443 662012 354509 662013
rect 354443 661948 354444 662012
rect 354508 661948 354509 662012
rect 354443 661947 354509 661948
rect 354446 655210 354506 661947
rect 354446 655150 354690 655210
rect 354630 654150 354690 655150
rect 354078 654090 354322 654150
rect 354262 345130 354322 654090
rect 354446 654090 354690 654150
rect 354446 644490 354506 654090
rect 354446 644430 354690 644490
rect 354630 644330 354690 644430
rect 354446 644270 354690 644330
rect 354446 635490 354506 644270
rect 354446 635430 354690 635490
rect 354630 634830 354690 635430
rect 354446 634770 354690 634830
rect 354446 625170 354506 634770
rect 354446 625110 354690 625170
rect 354630 624610 354690 625110
rect 354446 624550 354690 624610
rect 354446 615770 354506 624550
rect 354446 615710 354690 615770
rect 354630 615510 354690 615710
rect 354446 615450 354690 615510
rect 354446 605850 354506 615450
rect 354446 605790 354690 605850
rect 354630 605570 354690 605790
rect 354446 605510 354690 605570
rect 354446 596730 354506 605510
rect 354446 596670 354690 596730
rect 354630 596190 354690 596670
rect 354446 596130 354690 596190
rect 354446 586530 354506 596130
rect 354446 586470 354690 586530
rect 354630 585850 354690 586470
rect 354446 585790 354690 585850
rect 354446 577010 354506 585790
rect 354446 576950 354690 577010
rect 354630 576870 354690 576950
rect 354446 576810 354690 576870
rect 354446 567210 354506 576810
rect 354446 567150 354690 567210
rect 354630 566810 354690 567150
rect 354446 566750 354690 566810
rect 354446 557970 354506 566750
rect 354446 557910 354690 557970
rect 354630 557550 354690 557910
rect 354446 557490 354690 557550
rect 354446 547890 354506 557490
rect 354446 547830 354690 547890
rect 354630 547770 354690 547830
rect 354446 547710 354690 547770
rect 354446 538930 354506 547710
rect 354446 538870 354690 538930
rect 354630 538230 354690 538870
rect 354446 538170 354690 538230
rect 354446 528570 354506 538170
rect 354446 528510 354690 528570
rect 354630 528050 354690 528510
rect 354446 527990 354690 528050
rect 354446 519210 354506 527990
rect 354446 519150 354690 519210
rect 354630 518910 354690 519150
rect 354446 518850 354690 518910
rect 354446 509250 354506 518850
rect 354446 509190 354690 509250
rect 354630 509010 354690 509190
rect 354446 508950 354690 509010
rect 354446 500170 354506 508950
rect 354446 500110 354690 500170
rect 354630 499590 354690 500110
rect 354446 499530 354690 499590
rect 354446 489930 354506 499530
rect 354446 489870 354690 489930
rect 354630 489290 354690 489870
rect 354446 489230 354690 489290
rect 354446 480450 354506 489230
rect 354446 480390 354690 480450
rect 354630 480270 354690 480390
rect 354446 480210 354690 480270
rect 354446 470610 354506 480210
rect 354446 470550 354690 470610
rect 354630 470250 354690 470550
rect 354446 470190 354690 470250
rect 354446 461410 354506 470190
rect 354446 461350 354690 461410
rect 354630 460950 354690 461350
rect 354446 460890 354690 460950
rect 354446 451290 354506 460890
rect 354446 451230 354690 451290
rect 354630 450530 354690 451230
rect 354446 450470 354690 450530
rect 354446 442370 354506 450470
rect 354446 442310 354690 442370
rect 354630 441630 354690 442310
rect 354446 441570 354690 441630
rect 354446 431970 354506 441570
rect 354446 431910 354690 431970
rect 354630 431490 354690 431910
rect 354446 431430 354690 431490
rect 354446 422650 354506 431430
rect 354446 422590 354690 422650
rect 354630 422310 354690 422590
rect 354446 422250 354690 422310
rect 354446 412650 354506 422250
rect 354446 412590 354690 412650
rect 354630 412450 354690 412590
rect 354446 412390 354690 412450
rect 354446 403610 354506 412390
rect 354446 403550 354690 403610
rect 354630 402990 354690 403550
rect 354446 402930 354690 402990
rect 354446 393330 354506 402930
rect 354446 393270 354690 393330
rect 354630 392730 354690 393270
rect 354446 392670 354690 392730
rect 354446 383890 354506 392670
rect 354446 383830 354690 383890
rect 354630 383670 354690 383830
rect 354446 383610 354690 383670
rect 354446 374010 354506 383610
rect 354446 373950 354690 374010
rect 354630 373690 354690 373950
rect 354446 373630 354690 373690
rect 354446 364850 354506 373630
rect 354446 364790 354690 364850
rect 354630 364350 354690 364790
rect 354446 364290 354690 364350
rect 354446 354690 354506 364290
rect 354446 354630 354690 354690
rect 354630 353970 354690 354630
rect 354446 353910 354690 353970
rect 354446 345810 354506 353910
rect 354446 345750 354690 345810
rect 354262 345070 354506 345130
rect 354446 344450 354506 345070
rect 354262 344390 354506 344450
rect 354262 45930 354322 344390
rect 354630 343770 354690 345750
rect 354446 343710 354690 343770
rect 354446 335370 354506 343710
rect 354446 335310 354690 335370
rect 354630 334930 354690 335310
rect 354446 334870 354690 334930
rect 354446 326090 354506 334870
rect 354446 326030 354690 326090
rect 354630 325710 354690 326030
rect 354446 325650 354690 325710
rect 354446 316050 354506 325650
rect 354446 315990 354690 316050
rect 354630 315890 354690 315990
rect 354446 315830 354690 315890
rect 354446 307050 354506 315830
rect 354446 306990 354690 307050
rect 354630 306390 354690 306990
rect 354446 306330 354690 306390
rect 354446 296730 354506 306330
rect 354446 296670 354690 296730
rect 354630 296170 354690 296670
rect 354446 296110 354690 296170
rect 354446 287330 354506 296110
rect 354446 287270 354690 287330
rect 354630 287070 354690 287270
rect 354446 287010 354690 287070
rect 354446 277410 354506 287010
rect 354446 277350 354690 277410
rect 354630 277130 354690 277350
rect 354446 277070 354690 277130
rect 354446 268290 354506 277070
rect 354446 268230 354690 268290
rect 354630 267750 354690 268230
rect 354446 267690 354690 267750
rect 354446 258090 354506 267690
rect 354446 258030 354690 258090
rect 354630 257410 354690 258030
rect 354446 257350 354690 257410
rect 354446 248570 354506 257350
rect 354446 248510 354690 248570
rect 354630 248430 354690 248510
rect 354446 248370 354690 248430
rect 354446 238770 354506 248370
rect 354446 238710 354690 238770
rect 354630 238370 354690 238710
rect 354446 238310 354690 238370
rect 354446 229530 354506 238310
rect 354446 229470 354690 229530
rect 354630 229110 354690 229470
rect 354446 229050 354690 229110
rect 354446 219450 354506 229050
rect 354446 219390 354690 219450
rect 354630 219330 354690 219390
rect 354446 219270 354690 219330
rect 354446 210490 354506 219270
rect 354446 210430 354690 210490
rect 354630 209790 354690 210430
rect 354446 209730 354690 209790
rect 354446 200130 354506 209730
rect 354446 200070 354690 200130
rect 354630 199610 354690 200070
rect 354446 199550 354690 199610
rect 354446 190770 354506 199550
rect 354446 190710 354690 190770
rect 354630 190470 354690 190710
rect 354446 190410 354690 190470
rect 354446 180810 354506 190410
rect 354446 180750 354690 180810
rect 354630 180570 354690 180750
rect 354446 180510 354690 180570
rect 354446 171730 354506 180510
rect 354446 171670 354690 171730
rect 354630 171150 354690 171670
rect 354446 171090 354690 171150
rect 354446 161490 354506 171090
rect 354446 161430 354690 161490
rect 354630 160850 354690 161430
rect 354446 160790 354690 160850
rect 354446 152010 354506 160790
rect 354446 151950 354690 152010
rect 354630 151830 354690 151950
rect 354446 151770 354690 151830
rect 354446 142170 354506 151770
rect 354446 142110 354690 142170
rect 354630 141810 354690 142110
rect 354446 141750 354690 141810
rect 354446 132970 354506 141750
rect 354446 132910 354690 132970
rect 354630 132510 354690 132910
rect 354446 132450 354690 132510
rect 354446 122850 354506 132450
rect 354446 122790 354690 122850
rect 354630 122090 354690 122790
rect 354446 122030 354690 122090
rect 354446 113930 354506 122030
rect 354446 113870 354690 113930
rect 354630 113190 354690 113870
rect 354446 113130 354690 113190
rect 354446 103530 354506 113130
rect 354446 103470 354690 103530
rect 354630 103050 354690 103470
rect 354446 102990 354690 103050
rect 354446 94210 354506 102990
rect 354446 94150 354690 94210
rect 354630 93870 354690 94150
rect 354446 93810 354690 93870
rect 354446 84210 354506 93810
rect 354446 84150 354690 84210
rect 354630 84010 354690 84150
rect 354446 83950 354690 84010
rect 354446 75170 354506 83950
rect 354446 75110 354690 75170
rect 354630 74550 354690 75110
rect 354446 74490 354690 74550
rect 354446 64890 354506 74490
rect 354446 64830 354690 64890
rect 354630 64290 354690 64830
rect 354446 64230 354690 64290
rect 354446 55450 354506 64230
rect 354446 55390 354690 55450
rect 354630 55230 354690 55390
rect 354446 55170 354690 55230
rect 354446 51090 354506 55170
rect 354446 51030 354690 51090
rect 354262 45870 354506 45930
rect 354259 41444 354325 41445
rect 354259 41380 354260 41444
rect 354324 41380 354325 41444
rect 354259 41379 354325 41380
rect 353523 39132 353589 39133
rect 353523 39068 353524 39132
rect 353588 39068 353589 39132
rect 353523 39067 353589 39068
rect 354262 36005 354322 41379
rect 354259 36004 354325 36005
rect 354259 35940 354260 36004
rect 354324 35940 354325 36004
rect 354259 35939 354325 35940
rect 295931 33556 295997 33557
rect 295931 33492 295932 33556
rect 295996 33492 295997 33556
rect 295931 33491 295997 33492
rect 207611 8940 207677 8941
rect 207611 8876 207612 8940
rect 207676 8876 207677 8940
rect 207611 8875 207677 8876
rect 354446 6930 354506 45870
rect 354630 41445 354690 51030
rect 354814 43893 354874 663715
rect 355363 662420 355429 662421
rect 355363 662356 355364 662420
rect 355428 662356 355429 662420
rect 355363 662355 355429 662356
rect 355366 644490 355426 662355
rect 356099 662284 356165 662285
rect 356099 662220 356100 662284
rect 356164 662220 356165 662284
rect 356099 662219 356165 662220
rect 354998 644430 355426 644490
rect 354998 345030 355058 644430
rect 354998 344970 355426 345030
rect 355366 339690 355426 344970
rect 354998 339630 355426 339690
rect 354998 55230 355058 339630
rect 354998 55170 355242 55230
rect 354811 43892 354877 43893
rect 354811 43828 354812 43892
rect 354876 43828 354877 43892
rect 354811 43827 354877 43828
rect 355182 43349 355242 55170
rect 355179 43348 355245 43349
rect 355179 43284 355180 43348
rect 355244 43284 355245 43348
rect 355179 43283 355245 43284
rect 354627 41444 354693 41445
rect 354627 41380 354628 41444
rect 354692 41380 354693 41444
rect 354627 41379 354693 41380
rect 356102 40357 356162 662219
rect 358675 662148 358741 662149
rect 358675 662084 358676 662148
rect 358740 662084 358741 662148
rect 358675 662083 358741 662084
rect 356651 661876 356717 661877
rect 356651 661812 356652 661876
rect 356716 661812 356717 661876
rect 356651 661811 356717 661812
rect 356099 40356 356165 40357
rect 356099 40292 356100 40356
rect 356164 40292 356165 40356
rect 356099 40291 356165 40292
rect 354627 36004 354693 36005
rect 354627 35940 354628 36004
rect 354692 35940 354693 36004
rect 354627 35939 354693 35940
rect 354630 35733 354690 35939
rect 354627 35732 354693 35733
rect 354627 35668 354628 35732
rect 354692 35668 354693 35732
rect 354627 35667 354693 35668
rect 354627 26348 354693 26349
rect 354627 26284 354628 26348
rect 354692 26284 354693 26348
rect 354627 26283 354693 26284
rect 354630 26213 354690 26283
rect 354627 26212 354693 26213
rect 354627 26148 354628 26212
rect 354692 26148 354693 26212
rect 354627 26147 354693 26148
rect 354811 16692 354877 16693
rect 354811 16690 354812 16692
rect 354630 16630 354812 16690
rect 354630 16557 354690 16630
rect 354811 16628 354812 16630
rect 354876 16628 354877 16692
rect 354811 16627 354877 16628
rect 354627 16556 354693 16557
rect 354627 16492 354628 16556
rect 354692 16492 354693 16556
rect 354627 16491 354693 16492
rect 354627 7172 354693 7173
rect 354627 7108 354628 7172
rect 354692 7108 354693 7172
rect 354627 7107 354693 7108
rect 354262 6870 354506 6930
rect 55075 3908 55141 3909
rect 55075 3844 55076 3908
rect 55140 3844 55141 3908
rect 55075 3843 55141 3844
rect 42563 3500 42629 3501
rect 42563 3436 42564 3500
rect 42628 3436 42629 3500
rect 42563 3435 42629 3436
rect 39251 3364 39317 3365
rect 39251 3300 39252 3364
rect 39316 3300 39317 3364
rect 39251 3299 39317 3300
rect 354262 3229 354322 6870
rect 354630 6490 354690 7107
rect 354446 6430 354690 6490
rect 354446 5405 354506 6430
rect 354443 5404 354509 5405
rect 354443 5340 354444 5404
rect 354508 5340 354509 5404
rect 354443 5339 354509 5340
rect 354259 3228 354325 3229
rect 354259 3164 354260 3228
rect 354324 3164 354325 3228
rect 354259 3163 354325 3164
rect 356654 3093 356714 661811
rect 358678 39405 358738 662083
rect 358859 662012 358925 662013
rect 358859 661948 358860 662012
rect 358924 661948 358925 662012
rect 358859 661947 358925 661948
rect 358675 39404 358741 39405
rect 358675 39340 358676 39404
rect 358740 39340 358741 39404
rect 358675 39339 358741 39340
rect 358862 3909 358922 661947
rect 358859 3908 358925 3909
rect 358859 3844 358860 3908
rect 358924 3844 358925 3908
rect 358859 3843 358925 3844
rect 356651 3092 356717 3093
rect 356651 3028 356652 3092
rect 356716 3028 356717 3092
rect 356651 3027 356717 3028
rect 360702 2957 360762 664259
rect 362174 38861 362234 700027
rect 364931 699956 364997 699957
rect 364931 699892 364932 699956
rect 364996 699892 364997 699956
rect 364931 699891 364997 699892
rect 367691 699956 367757 699957
rect 367691 699892 367692 699956
rect 367756 699892 367757 699956
rect 367691 699891 367757 699892
rect 363459 664596 363525 664597
rect 363459 664532 363460 664596
rect 363524 664532 363525 664596
rect 363459 664531 363525 664532
rect 362171 38860 362237 38861
rect 362171 38796 362172 38860
rect 362236 38796 362237 38860
rect 362171 38795 362237 38796
rect 363462 3093 363522 664531
rect 364934 38725 364994 699891
rect 365667 699820 365733 699821
rect 365667 699756 365668 699820
rect 365732 699756 365733 699820
rect 365667 699755 365733 699756
rect 365670 39269 365730 699755
rect 366035 661876 366101 661877
rect 366035 661812 366036 661876
rect 366100 661812 366101 661876
rect 366035 661811 366101 661812
rect 366038 661197 366098 661811
rect 366035 661196 366101 661197
rect 366035 661132 366036 661196
rect 366100 661132 366101 661196
rect 366035 661131 366101 661132
rect 365667 39268 365733 39269
rect 365667 39204 365668 39268
rect 365732 39204 365733 39268
rect 365667 39203 365733 39204
rect 367694 39133 367754 699891
rect 368979 664732 369045 664733
rect 368979 664668 368980 664732
rect 369044 664668 369045 664732
rect 368979 664667 369045 664668
rect 367691 39132 367757 39133
rect 367691 39068 367692 39132
rect 367756 39068 367757 39132
rect 367691 39067 367757 39068
rect 364931 38724 364997 38725
rect 364931 38660 364932 38724
rect 364996 38660 364997 38724
rect 364931 38659 364997 38660
rect 368982 3909 369042 664667
rect 370454 42397 370514 700163
rect 402835 664324 402901 664325
rect 402835 664260 402836 664324
rect 402900 664260 402901 664324
rect 402835 664259 402901 664260
rect 394739 661876 394805 661877
rect 394739 661812 394740 661876
rect 394804 661812 394805 661876
rect 394739 661811 394805 661812
rect 370451 42396 370517 42397
rect 370451 42332 370452 42396
rect 370516 42332 370517 42396
rect 370451 42331 370517 42332
rect 394742 5541 394802 661811
rect 394739 5540 394805 5541
rect 394739 5476 394740 5540
rect 394804 5476 394805 5540
rect 394739 5475 394805 5476
rect 368979 3908 369045 3909
rect 368979 3844 368980 3908
rect 369044 3844 369045 3908
rect 368979 3843 369045 3844
rect 363459 3092 363525 3093
rect 363459 3028 363460 3092
rect 363524 3028 363525 3092
rect 363459 3027 363525 3028
rect 402838 2957 402898 664259
rect 405598 42397 405658 700843
rect 415899 700228 415965 700229
rect 415899 700164 415900 700228
rect 415964 700164 415965 700228
rect 415899 700163 415965 700164
rect 405595 42396 405661 42397
rect 405595 42332 405596 42396
rect 405660 42332 405661 42396
rect 405595 42331 405661 42332
rect 415902 40085 415962 700163
rect 467787 699820 467853 699821
rect 467787 699756 467788 699820
rect 467852 699756 467853 699820
rect 467787 699755 467853 699756
rect 488579 699820 488645 699821
rect 488579 699756 488580 699820
rect 488644 699756 488645 699820
rect 488579 699755 488645 699756
rect 436691 664460 436757 664461
rect 436691 664396 436692 664460
rect 436756 664396 436757 664460
rect 436691 664395 436757 664396
rect 425099 660380 425165 660381
rect 425099 660316 425100 660380
rect 425164 660316 425165 660380
rect 425099 660315 425165 660316
rect 415899 40084 415965 40085
rect 415899 40020 415900 40084
rect 415964 40020 415965 40084
rect 415899 40019 415965 40020
rect 425102 3093 425162 660315
rect 425099 3092 425165 3093
rect 425099 3028 425100 3092
rect 425164 3028 425165 3092
rect 425099 3027 425165 3028
rect 436694 2957 436754 664395
rect 443499 663916 443565 663917
rect 443499 663852 443500 663916
rect 443564 663852 443565 663916
rect 443499 663851 443565 663852
rect 440187 661876 440253 661877
rect 440187 661812 440188 661876
rect 440252 661812 440253 661876
rect 440187 661811 440253 661812
rect 440190 3093 440250 661811
rect 443502 6493 443562 663851
rect 451043 661876 451109 661877
rect 451043 661812 451044 661876
rect 451108 661812 451109 661876
rect 451043 661811 451109 661812
rect 460979 661876 461045 661877
rect 460979 661812 460980 661876
rect 461044 661812 461045 661876
rect 460979 661811 461045 661812
rect 466499 661876 466565 661877
rect 466499 661812 466500 661876
rect 466564 661812 466565 661876
rect 466499 661811 466565 661812
rect 443499 6492 443565 6493
rect 443499 6428 443500 6492
rect 443564 6428 443565 6492
rect 443499 6427 443565 6428
rect 451046 3773 451106 661811
rect 451043 3772 451109 3773
rect 451043 3708 451044 3772
rect 451108 3708 451109 3772
rect 451043 3707 451109 3708
rect 460982 3637 461042 661811
rect 466502 4045 466562 661811
rect 467790 39541 467850 699755
rect 488582 39813 488642 699755
rect 541019 663916 541085 663917
rect 541019 663852 541020 663916
rect 541084 663852 541085 663916
rect 541019 663851 541085 663852
rect 512131 661740 512197 661741
rect 512131 661676 512132 661740
rect 512196 661676 512197 661740
rect 512131 661675 512197 661676
rect 515259 661740 515325 661741
rect 515259 661676 515260 661740
rect 515324 661676 515325 661740
rect 515259 661675 515325 661676
rect 524459 661740 524525 661741
rect 524459 661676 524460 661740
rect 524524 661676 524525 661740
rect 524459 661675 524525 661676
rect 488579 39812 488645 39813
rect 488579 39748 488580 39812
rect 488644 39748 488645 39812
rect 488579 39747 488645 39748
rect 467787 39540 467853 39541
rect 467787 39476 467788 39540
rect 467852 39476 467853 39540
rect 467787 39475 467853 39476
rect 512134 4997 512194 661675
rect 512131 4996 512197 4997
rect 512131 4932 512132 4996
rect 512196 4932 512197 4996
rect 512131 4931 512197 4932
rect 466499 4044 466565 4045
rect 466499 3980 466500 4044
rect 466564 3980 466565 4044
rect 466499 3979 466565 3980
rect 515262 3637 515322 661675
rect 524462 5269 524522 661675
rect 541022 6357 541082 663851
rect 541755 661332 541821 661333
rect 541755 661268 541756 661332
rect 541820 661268 541821 661332
rect 541755 661267 541821 661268
rect 541758 473370 541818 661267
rect 541574 473310 541818 473370
rect 541574 468890 541634 473310
rect 541942 471885 542002 700979
rect 542859 700636 542925 700637
rect 542859 700572 542860 700636
rect 542924 700572 542925 700636
rect 542859 700571 542925 700572
rect 542491 700500 542557 700501
rect 542491 700436 542492 700500
rect 542556 700436 542557 700500
rect 542491 700435 542557 700436
rect 542123 660244 542189 660245
rect 542123 660180 542124 660244
rect 542188 660180 542189 660244
rect 542123 660179 542189 660180
rect 542307 660244 542373 660245
rect 542307 660180 542308 660244
rect 542372 660180 542373 660244
rect 542307 660179 542373 660180
rect 542126 653445 542186 660179
rect 542123 653444 542189 653445
rect 542123 653380 542124 653444
rect 542188 653380 542189 653444
rect 542123 653379 542189 653380
rect 542310 592925 542370 660179
rect 542307 592924 542373 592925
rect 542307 592860 542308 592924
rect 542372 592860 542373 592924
rect 542307 592859 542373 592860
rect 542307 587756 542373 587757
rect 542307 587692 542308 587756
rect 542372 587692 542373 587756
rect 542307 587691 542373 587692
rect 542123 482220 542189 482221
rect 542123 482156 542124 482220
rect 542188 482156 542189 482220
rect 542123 482155 542189 482156
rect 541939 471884 542005 471885
rect 541939 471820 541940 471884
rect 542004 471820 542005 471884
rect 541939 471819 542005 471820
rect 541574 468830 541818 468890
rect 541758 468349 541818 468830
rect 541755 468348 541821 468349
rect 541755 468284 541756 468348
rect 541820 468284 541821 468348
rect 541755 468283 541821 468284
rect 542126 468210 542186 482155
rect 541574 468150 542186 468210
rect 541574 443010 541634 468150
rect 541755 468076 541821 468077
rect 541755 468012 541756 468076
rect 541820 468012 541821 468076
rect 541755 468011 541821 468012
rect 541758 445090 541818 468011
rect 541939 466308 542005 466309
rect 541939 466244 541940 466308
rect 542004 466244 542005 466308
rect 541939 466243 542005 466244
rect 541942 445773 542002 466243
rect 541939 445772 542005 445773
rect 541939 445708 541940 445772
rect 542004 445708 542005 445772
rect 541939 445707 542005 445708
rect 541758 445030 542002 445090
rect 541755 444412 541821 444413
rect 541755 444348 541756 444412
rect 541820 444348 541821 444412
rect 541755 444347 541821 444348
rect 541206 442950 541634 443010
rect 541206 440330 541266 442950
rect 541758 442509 541818 444347
rect 541755 442508 541821 442509
rect 541755 442444 541756 442508
rect 541820 442444 541821 442508
rect 541755 442443 541821 442444
rect 541206 440270 541818 440330
rect 541758 439109 541818 440270
rect 541755 439108 541821 439109
rect 541755 439044 541756 439108
rect 541820 439044 541821 439108
rect 541755 439043 541821 439044
rect 541755 438972 541821 438973
rect 541755 438970 541756 438972
rect 541206 438910 541756 438970
rect 541019 6356 541085 6357
rect 541019 6292 541020 6356
rect 541084 6292 541085 6356
rect 541019 6291 541085 6292
rect 541206 6221 541266 438910
rect 541755 438908 541756 438910
rect 541820 438908 541821 438972
rect 541755 438907 541821 438908
rect 541755 438156 541821 438157
rect 541755 438092 541756 438156
rect 541820 438092 541821 438156
rect 541755 438091 541821 438092
rect 541758 433350 541818 438091
rect 541574 433290 541818 433350
rect 541942 433350 542002 445030
rect 541942 433290 542186 433350
rect 541574 44301 541634 433290
rect 542126 431970 542186 433290
rect 541758 431910 542186 431970
rect 541758 291141 541818 431910
rect 541755 291140 541821 291141
rect 541755 291076 541756 291140
rect 541820 291076 541821 291140
rect 541755 291075 541821 291076
rect 541755 150516 541821 150517
rect 541755 150452 541756 150516
rect 541820 150452 541821 150516
rect 541755 150451 541821 150452
rect 541758 44437 541818 150451
rect 541939 49604 542005 49605
rect 541939 49540 541940 49604
rect 542004 49540 542005 49604
rect 541939 49539 542005 49540
rect 541755 44436 541821 44437
rect 541755 44372 541756 44436
rect 541820 44372 541821 44436
rect 541755 44371 541821 44372
rect 541571 44300 541637 44301
rect 541571 44236 541572 44300
rect 541636 44236 541637 44300
rect 541571 44235 541637 44236
rect 541942 44029 542002 49539
rect 541939 44028 542005 44029
rect 541939 43964 541940 44028
rect 542004 43964 542005 44028
rect 541939 43963 542005 43964
rect 542310 10301 542370 587691
rect 542494 284205 542554 700435
rect 542675 296716 542741 296717
rect 542675 296652 542676 296716
rect 542740 296652 542741 296716
rect 542675 296651 542741 296652
rect 542491 284204 542557 284205
rect 542491 284140 542492 284204
rect 542556 284140 542557 284204
rect 542491 284139 542557 284140
rect 542678 44573 542738 296651
rect 542862 139501 542922 700571
rect 543779 699820 543845 699821
rect 543779 699756 543780 699820
rect 543844 699756 543845 699820
rect 543779 699755 543845 699756
rect 543595 660516 543661 660517
rect 543595 660452 543596 660516
rect 543660 660452 543661 660516
rect 543595 660451 543661 660452
rect 543043 369204 543109 369205
rect 543043 369140 543044 369204
rect 543108 369140 543109 369204
rect 543043 369139 543109 369140
rect 542859 139500 542925 139501
rect 542859 139436 542860 139500
rect 542924 139436 542925 139500
rect 542859 139435 542925 139436
rect 542675 44572 542741 44573
rect 542675 44508 542676 44572
rect 542740 44508 542741 44572
rect 542675 44507 542741 44508
rect 542307 10300 542373 10301
rect 542307 10236 542308 10300
rect 542372 10236 542373 10300
rect 542307 10235 542373 10236
rect 541203 6220 541269 6221
rect 541203 6156 541204 6220
rect 541268 6156 541269 6220
rect 541203 6155 541269 6156
rect 524459 5268 524525 5269
rect 524459 5204 524460 5268
rect 524524 5204 524525 5268
rect 524459 5203 524525 5204
rect 460979 3636 461045 3637
rect 460979 3572 460980 3636
rect 461044 3572 461045 3636
rect 460979 3571 461045 3572
rect 515259 3636 515325 3637
rect 515259 3572 515260 3636
rect 515324 3572 515325 3636
rect 515259 3571 515325 3572
rect 543046 3501 543106 369139
rect 543598 191725 543658 660451
rect 543595 191724 543661 191725
rect 543595 191660 543596 191724
rect 543660 191660 543661 191724
rect 543595 191659 543661 191660
rect 543782 42125 543842 699755
rect 545067 664188 545133 664189
rect 545067 664124 545068 664188
rect 545132 664124 545133 664188
rect 545067 664123 545133 664124
rect 544331 660924 544397 660925
rect 544331 660860 544332 660924
rect 544396 660860 544397 660924
rect 544331 660859 544397 660860
rect 543963 543012 544029 543013
rect 543963 542948 543964 543012
rect 544028 542948 544029 543012
rect 543963 542947 544029 542948
rect 543779 42124 543845 42125
rect 543779 42060 543780 42124
rect 543844 42060 543845 42124
rect 543779 42059 543845 42060
rect 543966 4861 544026 542947
rect 544147 471476 544213 471477
rect 544147 471412 544148 471476
rect 544212 471412 544213 471476
rect 544147 471411 544213 471412
rect 544150 43485 544210 471411
rect 544334 234157 544394 660859
rect 544515 660380 544581 660381
rect 544515 660316 544516 660380
rect 544580 660316 544581 660380
rect 544515 660315 544581 660316
rect 544518 261085 544578 660315
rect 544515 261084 544581 261085
rect 544515 261020 544516 261084
rect 544580 261020 544581 261084
rect 544515 261019 544581 261020
rect 544331 234156 544397 234157
rect 544331 234092 544332 234156
rect 544396 234092 544397 234156
rect 544331 234091 544397 234092
rect 544331 135556 544397 135557
rect 544331 135492 544332 135556
rect 544396 135492 544397 135556
rect 544331 135491 544397 135492
rect 544334 49605 544394 135491
rect 544331 49604 544397 49605
rect 544331 49540 544332 49604
rect 544396 49540 544397 49604
rect 544331 49539 544397 49540
rect 544147 43484 544213 43485
rect 544147 43420 544148 43484
rect 544212 43420 544213 43484
rect 544147 43419 544213 43420
rect 545070 33829 545130 664123
rect 545619 661060 545685 661061
rect 545619 660996 545620 661060
rect 545684 660996 545685 661060
rect 545619 660995 545685 660996
rect 545251 583268 545317 583269
rect 545251 583204 545252 583268
rect 545316 583204 545317 583268
rect 545251 583203 545317 583204
rect 545067 33828 545133 33829
rect 545067 33764 545068 33828
rect 545132 33764 545133 33828
rect 545067 33763 545133 33764
rect 545254 5133 545314 583203
rect 545622 16693 545682 660995
rect 545619 16692 545685 16693
rect 545619 16628 545620 16692
rect 545684 16628 545685 16692
rect 545619 16627 545685 16628
rect 545251 5132 545317 5133
rect 545251 5068 545252 5132
rect 545316 5068 545317 5132
rect 545251 5067 545317 5068
rect 543963 4860 544029 4861
rect 543963 4796 543964 4860
rect 544028 4796 544029 4860
rect 543963 4795 544029 4796
rect 543043 3500 543109 3501
rect 543043 3436 543044 3500
rect 543108 3436 543109 3500
rect 543043 3435 543109 3436
rect 440187 3092 440253 3093
rect 440187 3028 440188 3092
rect 440252 3028 440253 3092
rect 440187 3027 440253 3028
rect 360699 2956 360765 2957
rect 360699 2892 360700 2956
rect 360764 2892 360765 2956
rect 360699 2891 360765 2892
rect 402835 2956 402901 2957
rect 402835 2892 402836 2956
rect 402900 2892 402901 2956
rect 402835 2891 402901 2892
rect 436691 2956 436757 2957
rect 436691 2892 436692 2956
rect 436756 2892 436757 2956
rect 436691 2891 436757 2892
use top  TopSoC
timestamp 1633664140
transform 1 0 42000 0 1 42000
box -960 -960 500960 620960
<< labels >>
rlabel metal2 s 405894 703520 406006 704960 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 647036 584960 647276 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 224076 584960 224316 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 139646 -960 139758 480 8 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 422638 -960 422750 480 8 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 445822 703520 445934 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal3 s 583520 76380 584960 76620 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 109838 -960 109950 480 8 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 66414 -960 66526 480 8 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 545734 -960 545846 480 8 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s 583520 568428 584960 568668 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal2 s 359158 703520 359270 704960 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 152268 480 152508 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s 583520 145196 584960 145436 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 409206 703520 409318 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 172950 -960 173062 480 8 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal2 s 525678 703520 525790 704960 6 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal2 s 212878 -960 212990 480 8 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s 583520 627452 584960 627692 6 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s 583520 701164 584960 701404 6 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal2 s 13054 703520 13166 704960 6 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal2 s 232750 703520 232862 704960 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s -960 526268 480 526508 4 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal2 s 296046 703520 296158 704960 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s -960 619836 480 620076 4 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s -960 536060 480 536300 4 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 91068 584960 91308 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal3 s -960 98140 480 98380 4 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 563532 584960 563772 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 583116 584960 583356 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s -960 48908 480 49148 4 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 238764 584960 239004 6 io_in[11]
port 31 nsew signal input
rlabel metal2 s 472318 703520 472430 704960 6 io_in[12]
port 32 nsew signal input
rlabel metal2 s 192822 703520 192934 704960 6 io_in[13]
port 33 nsew signal input
rlabel metal2 s 199446 703520 199558 704960 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 86286 703520 86398 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 19678 703520 19790 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 219502 703520 219614 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal3 s -960 551020 480 551260 4 io_in[18]
port 38 nsew signal input
rlabel metal2 s 222814 703520 222926 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal2 s 66230 703520 66342 704960 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 359342 -960 359454 480 8 io_in[20]
port 41 nsew signal input
rlabel metal3 s 583520 533884 584960 534124 6 io_in[21]
port 42 nsew signal input
rlabel metal3 s 583520 105756 584960 105996 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 193006 -960 193118 480 8 io_in[23]
port 44 nsew signal input
rlabel metal2 s 309294 703520 309406 704960 6 io_in[24]
port 45 nsew signal input
rlabel metal3 s 583520 17356 584960 17596 6 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 9740 480 9980 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 413116 480 413356 4 io_in[27]
port 48 nsew signal input
rlabel metal2 s 568918 703520 569030 704960 6 io_in[28]
port 49 nsew signal input
rlabel metal3 s 583520 81276 584960 81516 6 io_in[29]
port 50 nsew signal input
rlabel metal3 s -960 659276 480 659516 4 io_in[2]
port 51 nsew signal input
rlabel metal2 s 572230 703520 572342 704960 6 io_in[30]
port 52 nsew signal input
rlabel metal2 s 126214 703520 126326 704960 6 io_in[31]
port 53 nsew signal input
rlabel metal3 s 583520 140300 584960 140540 6 io_in[32]
port 54 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 io_in[33]
port 55 nsew signal input
rlabel metal2 s 43046 703520 43158 704960 6 io_in[34]
port 56 nsew signal input
rlabel metal2 s 412518 703520 412630 704960 6 io_in[35]
port 57 nsew signal input
rlabel metal2 s 245998 703520 246110 704960 6 io_in[36]
port 58 nsew signal input
rlabel metal3 s 583520 61692 584960 61932 6 io_in[37]
port 59 nsew signal input
rlabel metal2 s 512430 703520 512542 704960 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s -960 698444 480 698684 4 io_in[4]
port 61 nsew signal input
rlabel metal2 s 356030 -960 356142 480 8 io_in[5]
port 62 nsew signal input
rlabel metal3 s -960 363884 480 364124 4 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 696268 584960 696508 6 io_in[7]
port 64 nsew signal input
rlabel metal2 s 425950 -960 426062 480 8 io_in[8]
port 65 nsew signal input
rlabel metal2 s 409390 -960 409502 480 8 io_in[9]
port 66 nsew signal input
rlabel metal2 s 555670 703520 555782 704960 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal2 s 129710 -960 129822 480 8 io_oeb[10]
port 68 nsew signal tristate
rlabel metal2 s 99718 -960 99830 480 8 io_oeb[11]
port 69 nsew signal tristate
rlabel metal2 s 529174 -960 529286 480 8 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 292892 584960 293132 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 548844 584960 549084 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal3 s -960 546124 480 546364 4 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 442694 -960 442806 480 8 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 565790 -960 565902 480 8 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 96222 703520 96334 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 545550 703520 545662 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal2 s 3118 703520 3230 704960 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal3 s -960 24428 480 24668 4 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 302854 -960 302966 480 8 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 16550 -960 16662 480 8 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 334508 480 334748 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s 583520 514300 584960 514540 6 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 245836 480 246076 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s 583520 263244 584960 263484 6 io_oeb[27]
port 86 nsew signal tristate
rlabel metal2 s 136150 703520 136262 704960 6 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 206396 480 206636 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s -960 580396 480 580636 4 io_oeb[2]
port 89 nsew signal tristate
rlabel metal2 s 32926 703520 33038 704960 6 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s 583520 622556 584960 622796 6 io_oeb[31]
port 91 nsew signal tristate
rlabel metal2 s 532302 703520 532414 704960 6 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s 583520 36940 584960 37180 6 io_oeb[33]
port 93 nsew signal tristate
rlabel metal2 s 325854 703520 325966 704960 6 io_oeb[34]
port 94 nsew signal tristate
rlabel metal2 s 156206 703520 156318 704960 6 io_oeb[35]
port 95 nsew signal tristate
rlabel metal2 s 259614 -960 259726 480 8 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 703612 480 703852 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal2 s 79662 703520 79774 704960 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 573324 584960 573564 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal2 s 435702 703520 435814 704960 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s -960 565708 480 565948 4 io_oeb[6]
port 101 nsew signal tristate
rlabel metal2 s 239558 -960 239670 480 8 io_oeb[7]
port 102 nsew signal tristate
rlabel metal2 s 46542 -960 46654 480 8 io_oeb[8]
port 103 nsew signal tristate
rlabel metal2 s 515926 -960 516038 480 8 io_oeb[9]
port 104 nsew signal tristate
rlabel metal2 s 292734 703520 292846 704960 6 io_out[0]
port 105 nsew signal tristate
rlabel metal2 s 475998 -960 476110 480 8 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s -960 108204 480 108444 4 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s -960 511580 480 511820 4 io_out[12]
port 108 nsew signal tristate
rlabel metal2 s 49670 703520 49782 704960 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 479756 584960 479996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 475814 703520 475926 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 49854 -960 49966 480 8 io_out[16]
port 112 nsew signal tristate
rlabel metal3 s -960 457452 480 457692 4 io_out[17]
port 113 nsew signal tristate
rlabel metal3 s -960 250732 480 250972 4 io_out[18]
port 114 nsew signal tristate
rlabel metal3 s 583520 337228 584960 337468 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s -960 462348 480 462588 4 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 79846 -960 79958 480 8 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 99534 703520 99646 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 26486 -960 26598 480 8 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s 583520 474860 584960 475100 6 io_out[24]
port 121 nsew signal tristate
rlabel metal2 s 242686 703520 242798 704960 6 io_out[25]
port 122 nsew signal tristate
rlabel metal2 s 319230 703520 319342 704960 6 io_out[26]
port 123 nsew signal tristate
rlabel metal2 s 389334 -960 389446 480 8 io_out[27]
port 124 nsew signal tristate
rlabel metal2 s 209382 703520 209494 704960 6 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s 583520 71484 584960 71724 6 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 460172 584960 460412 6 io_out[2]
port 127 nsew signal tristate
rlabel metal2 s 69726 -960 69838 480 8 io_out[30]
port 128 nsew signal tristate
rlabel metal2 s 209566 -960 209678 480 8 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s 583520 445484 584960 445724 6 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s 583520 283100 584960 283340 6 io_out[33]
port 131 nsew signal tristate
rlabel metal2 s 376086 -960 376198 480 8 io_out[34]
port 132 nsew signal tristate
rlabel metal2 s 83158 -960 83270 480 8 io_out[35]
port 133 nsew signal tristate
rlabel metal2 s 482438 703520 482550 704960 6 io_out[36]
port 134 nsew signal tristate
rlabel metal2 s 136334 -960 136446 480 8 io_out[37]
port 135 nsew signal tristate
rlabel metal2 s 133022 -960 133134 480 8 io_out[3]
port 136 nsew signal tristate
rlabel metal2 s 33110 -960 33222 480 8 io_out[4]
port 137 nsew signal tristate
rlabel metal2 s 425766 703520 425878 704960 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s -960 236044 480 236284 4 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 420732 584960 420972 6 io_out[7]
port 140 nsew signal tristate
rlabel metal2 s 269550 -960 269662 480 8 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 179740 584960 179980 6 io_out[9]
port 142 nsew signal tristate
rlabel metal3 s -960 501788 480 502028 4 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 212694 703520 212806 704960 6 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 279302 703520 279414 704960 6 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 206070 703520 206182 704960 6 la_data_in[102]
port 146 nsew signal input
rlabel metal3 s 583520 657100 584960 657340 6 la_data_in[103]
port 147 nsew signal input
rlabel metal3 s 583520 248556 584960 248796 6 la_data_in[104]
port 148 nsew signal input
rlabel metal3 s -960 221356 480 221596 4 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 52982 703520 53094 704960 6 la_data_in[106]
port 150 nsew signal input
rlabel metal3 s -960 383740 480 383980 4 la_data_in[107]
port 151 nsew signal input
rlabel metal3 s -960 649484 480 649724 4 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 196134 703520 196246 704960 6 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 73038 703520 73150 704960 6 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 355846 703520 355958 704960 6 la_data_in[111]
port 156 nsew signal input
rlabel metal3 s -960 39116 480 39356 4 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 93094 -960 93206 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal3 s -960 531164 480 531404 4 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 342782 -960 342894 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal3 s 583520 666892 584960 667132 6 la_data_in[116]
port 161 nsew signal input
rlabel metal3 s 583520 268140 584960 268380 6 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 309478 -960 309590 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal3 s 583520 440588 584960 440828 6 la_data_in[119]
port 164 nsew signal input
rlabel metal3 s -960 427804 480 428044 4 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 269366 703520 269478 704960 6 la_data_in[120]
port 166 nsew signal input
rlabel metal3 s 583520 504508 584960 504748 6 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 252622 703520 252734 704960 6 la_data_in[122]
port 168 nsew signal input
rlabel metal3 s 583520 425628 584960 425868 6 la_data_in[123]
port 169 nsew signal input
rlabel metal3 s 583520 243660 584960 243900 6 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 382710 -960 382822 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 452446 703520 452558 704960 6 la_data_in[126]
port 172 nsew signal input
rlabel metal3 s 583520 12460 584960 12700 6 la_data_in[127]
port 173 nsew signal input
rlabel metal3 s -960 304860 480 305100 4 la_data_in[12]
port 174 nsew signal input
rlabel metal3 s 583520 450380 584960 450620 6 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 508934 703520 509046 704960 6 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 239374 703520 239486 704960 6 la_data_in[15]
port 177 nsew signal input
rlabel metal3 s 583520 528988 584960 529228 6 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 542422 -960 542534 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 535798 -960 535910 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 352534 703520 352646 704960 6 la_data_in[19]
port 181 nsew signal input
rlabel metal3 s -960 654380 480 654620 4 la_data_in[1]
port 182 nsew signal input
rlabel metal3 s -960 162332 480 162572 4 la_data_in[20]
port 183 nsew signal input
rlabel metal3 s 583520 22252 584960 22492 6 la_data_in[21]
port 184 nsew signal input
rlabel metal3 s -960 467244 480 467484 4 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 76350 703520 76462 704960 6 la_data_in[23]
port 186 nsew signal input
rlabel metal3 s -960 285276 480 285516 4 la_data_in[24]
port 187 nsew signal input
rlabel metal3 s -960 68764 480 69004 4 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 259430 703520 259542 704960 6 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 232934 -960 233046 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal3 s 583520 312476 584960 312716 6 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 162830 703520 162942 704960 6 la_data_in[29]
port 192 nsew signal input
rlabel metal3 s -960 226252 480 226492 4 la_data_in[2]
port 193 nsew signal input
rlabel metal3 s -960 142476 480 142716 4 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 199630 -960 199742 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 322542 703520 322654 704960 6 la_data_in[32]
port 196 nsew signal input
rlabel metal3 s -960 634524 480 634764 4 la_data_in[33]
port 197 nsew signal input
rlabel metal3 s -960 585292 480 585532 4 la_data_in[34]
port 198 nsew signal input
rlabel metal3 s 583520 159884 584960 160124 6 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 432574 -960 432686 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 246182 -960 246294 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 92910 703520 93022 704960 6 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 36422 703520 36534 704960 6 la_data_in[39]
port 203 nsew signal input
rlabel metal3 s 583520 327436 584960 327676 6 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 262742 703520 262854 704960 6 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 176078 703520 176190 704960 6 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal3 s 583520 189532 584960 189772 6 la_data_in[43]
port 208 nsew signal input
rlabel metal3 s -960 63868 480 64108 4 la_data_in[44]
port 209 nsew signal input
rlabel metal3 s 583520 361708 584960 361948 6 la_data_in[45]
port 210 nsew signal input
rlabel metal3 s -960 265420 480 265660 4 la_data_in[46]
port 211 nsew signal input
rlabel metal3 s 583520 386460 584960 386700 6 la_data_in[47]
port 212 nsew signal input
rlabel metal3 s -960 422908 480 423148 4 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 129526 703520 129638 704960 6 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 346094 -960 346206 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 575542 703520 575654 704960 6 la_data_in[50]
port 216 nsew signal input
rlabel metal3 s -960 506684 480 506924 4 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 39734 703520 39846 704960 6 la_data_in[52]
port 218 nsew signal input
rlabel metal3 s -960 83452 480 83692 4 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 3302 -960 3414 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal3 s 583520 435692 584960 435932 6 la_data_in[55]
port 221 nsew signal input
rlabel metal3 s -960 570604 480 570844 4 la_data_in[56]
port 222 nsew signal input
rlabel metal3 s 583520 617660 584960 617900 6 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 73222 -960 73334 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal3 s 583520 356812 584960 357052 6 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 379214 703520 379326 704960 6 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal3 s 583520 415836 584960 416076 6 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 509118 -960 509230 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal3 s 583520 322268 584960 322508 6 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 395774 703520 395886 704960 6 la_data_in[64]
port 231 nsew signal input
rlabel metal3 s -960 516476 480 516716 4 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 552358 703520 552470 704960 6 la_data_in[66]
port 233 nsew signal input
rlabel metal3 s -960 418012 480 418252 4 la_data_in[67]
port 234 nsew signal input
rlabel metal3 s -960 595356 480 595596 4 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 505806 -960 505918 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal3 s 583520 174844 584960 175084 6 la_data_in[6]
port 237 nsew signal input
rlabel metal3 s 583520 553740 584960 553980 6 la_data_in[70]
port 238 nsew signal input
rlabel metal3 s 583520 598076 584960 598316 6 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 459070 703520 459182 704960 6 la_data_in[72]
port 240 nsew signal input
rlabel metal3 s -960 78556 480 78796 4 la_data_in[73]
port 241 nsew signal input
rlabel metal3 s 583520 204220 584960 204460 6 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 202758 703520 202870 704960 6 la_data_in[75]
port 243 nsew signal input
rlabel metal3 s 583520 7564 584960 7804 6 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 505622 703520 505734 704960 6 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 286110 -960 286222 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal3 s 583520 538780 584960 539020 6 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 279486 -960 279598 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal3 s -960 93244 480 93484 4 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 525862 -960 525974 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal3 s 583520 228972 584960 229212 6 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 535614 703520 535726 704960 6 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 469190 -960 469302 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 236062 703520 236174 704960 6 la_data_in[85]
port 254 nsew signal input
rlabel metal3 s 583520 351916 584960 352156 6 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 449134 703520 449246 704960 6 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 216006 703520 216118 704960 6 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 382526 703520 382638 704960 6 la_data_in[89]
port 258 nsew signal input
rlabel metal3 s -960 398428 480 398668 4 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 459254 -960 459366 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal3 s -960 452556 480 452796 4 la_data_in[91]
port 261 nsew signal input
rlabel metal3 s 583520 519196 584960 519436 6 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 285926 703520 286038 704960 6 la_data_in[93]
port 263 nsew signal input
rlabel metal3 s -960 349196 480 349436 4 la_data_in[94]
port 264 nsew signal input
rlabel metal3 s 583520 637244 584960 637484 6 la_data_in[95]
port 265 nsew signal input
rlabel metal3 s -960 560812 480 561052 4 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 422454 703520 422566 704960 6 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 229622 -960 229734 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal3 s -960 610044 480 610284 4 la_data_in[99]
port 269 nsew signal input
rlabel metal3 s 583520 302684 584960 302924 6 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 372590 703520 372702 704960 6 la_data_out[0]
port 271 nsew signal tristate
rlabel metal3 s 583520 376396 584960 376636 6 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 189694 -960 189806 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 103030 -960 103142 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal3 s 583520 130508 584960 130748 6 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 519054 703520 519166 704960 6 la_data_out[104]
port 276 nsew signal tristate
rlabel metal3 s 583520 56796 584960 57036 6 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 126398 -960 126510 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal3 s 583520 287996 584960 288236 6 la_data_out[107]
port 279 nsew signal tristate
rlabel metal3 s 583520 430524 584960 430764 6 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 442510 703520 442622 704960 6 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 362654 -960 362766 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal3 s -960 329612 480 329852 4 la_data_out[110]
port 283 nsew signal tristate
rlabel metal3 s 583520 100860 584960 101100 6 la_data_out[111]
port 284 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 166326 -960 166438 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 89598 703520 89710 704960 6 la_data_out[114]
port 287 nsew signal tristate
rlabel metal3 s 583520 51628 584960 51868 6 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 336158 -960 336270 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 106158 703520 106270 704960 6 la_data_out[117]
port 290 nsew signal tristate
rlabel metal3 s 583520 297788 584960 298028 6 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 499182 -960 499294 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal3 s 583520 165052 584960 165292 6 la_data_out[11]
port 293 nsew signal tristate
rlabel metal3 s -960 177020 480 177260 4 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 216190 -960 216302 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal3 s -960 34220 480 34460 4 la_data_out[122]
port 296 nsew signal tristate
rlabel metal3 s 583520 632348 584960 632588 6 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 542238 703520 542350 704960 6 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 59606 703520 59718 704960 6 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 152894 703520 153006 704960 6 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 139462 703520 139574 704960 6 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 186382 -960 186494 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 512614 -960 512726 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 16366 703520 16478 704960 6 la_data_out[14]
port 304 nsew signal tristate
rlabel metal3 s -960 555916 480 556156 4 la_data_out[15]
port 305 nsew signal tristate
rlabel metal3 s 583520 396252 584960 396492 6 la_data_out[16]
port 306 nsew signal tristate
rlabel metal3 s 583520 342124 584960 342364 6 la_data_out[17]
port 307 nsew signal tristate
rlabel metal3 s -960 216460 480 216700 4 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 146270 703520 146382 704960 6 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 552542 -960 552654 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 339286 703520 339398 704960 6 la_data_out[20]
port 311 nsew signal tristate
rlabel metal3 s 583520 110924 584960 111164 6 la_data_out[21]
port 312 nsew signal tristate
rlabel metal3 s -960 639420 480 639660 4 la_data_out[22]
port 313 nsew signal tristate
rlabel metal3 s 583520 115820 584960 116060 6 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 492558 -960 492670 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 522366 703520 522478 704960 6 la_data_out[25]
port 316 nsew signal tristate
rlabel metal3 s -960 447660 480 447900 4 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 166142 703520 166254 704960 6 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 256302 -960 256414 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 252806 -960 252918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 395958 -960 396070 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 332662 703520 332774 704960 6 la_data_out[30]
port 322 nsew signal tristate
rlabel metal3 s -960 290172 480 290412 4 la_data_out[31]
port 323 nsew signal tristate
rlabel metal3 s -960 354092 480 354332 4 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 385838 703520 385950 704960 6 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 262926 -960 263038 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal3 s 583520 27148 584960 27388 6 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 132838 703520 132950 704960 6 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 489246 -960 489358 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 539110 -960 539222 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal3 s 583520 2668 584960 2908 6 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 249310 703520 249422 704960 6 la_data_out[3]
port 332 nsew signal tristate
rlabel metal3 s 583520 253452 584960 253692 6 la_data_out[40]
port 333 nsew signal tristate
rlabel metal3 s -960 113100 480 113340 4 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 69542 703520 69654 704960 6 la_data_out[42]
port 335 nsew signal tristate
rlabel metal3 s -960 73660 480 73900 4 la_data_out[43]
port 336 nsew signal tristate
rlabel metal3 s -960 393532 480 393772 4 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 312790 -960 312902 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 179390 703520 179502 704960 6 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 56478 -960 56590 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 335974 703520 336086 704960 6 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 46358 703520 46470 704960 6 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 528990 703520 529102 704960 6 la_data_out[4]
port 343 nsew signal tristate
rlabel metal3 s -960 295068 480 295308 4 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal3 s -960 103036 480 103276 4 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 419142 703520 419254 704960 6 la_data_out[53]
port 347 nsew signal tristate
rlabel metal3 s -960 487100 480 487340 4 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 169638 -960 169750 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 349406 -960 349518 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 256118 703520 256230 704960 6 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 122902 703520 123014 704960 6 la_data_out[58]
port 352 nsew signal tristate
rlabel metal3 s -960 388636 480 388876 4 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 296230 -960 296342 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 289422 -960 289534 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 502310 703520 502422 704960 6 la_data_out[61]
port 356 nsew signal tristate
rlabel metal3 s -960 147372 480 147612 4 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 485750 703520 485862 704960 6 la_data_out[63]
port 358 nsew signal tristate
rlabel metal3 s -960 496892 480 497132 4 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 435886 -960 435998 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 485934 -960 486046 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal3 s 583520 391356 584960 391596 6 la_data_out[67]
port 362 nsew signal tristate
rlabel metal3 s 583520 135404 584960 135644 6 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 172766 703520 172878 704960 6 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 266238 -960 266350 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 392646 -960 392758 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 202942 -960 203054 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 22990 703520 23102 704960 6 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 299542 -960 299654 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 416014 -960 416126 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 332846 -960 332958 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 146454 -960 146566 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 116278 703520 116390 704960 6 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 276174 -960 276286 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal3 s -960 122892 480 123132 4 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 522550 -960 522662 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal3 s 583520 125612 584960 125852 6 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 182886 703520 182998 704960 6 la_data_out[81]
port 378 nsew signal tristate
rlabel metal3 s -960 58972 480 59212 4 la_data_out[82]
port 379 nsew signal tristate
rlabel metal3 s -960 683756 480 683996 4 la_data_out[83]
port 380 nsew signal tristate
rlabel metal3 s -960 260524 480 260764 4 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 549046 703520 549158 704960 6 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 449318 -960 449430 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal3 s 583520 681580 584960 681820 6 la_data_out[87]
port 384 nsew signal tristate
rlabel metal3 s -960 137580 480 137820 4 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 549230 -960 549342 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal3 s 583520 371500 584960 371740 6 la_data_out[8]
port 387 nsew signal tristate
rlabel metal3 s -960 664172 480 664412 4 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 226126 703520 226238 704960 6 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 289238 703520 289350 704960 6 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 26302 703520 26414 704960 6 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 412702 -960 412814 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 465878 -960 465990 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 315918 703520 316030 704960 6 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 159702 -960 159814 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 578854 703520 578966 704960 6 la_data_out[98]
port 396 nsew signal tristate
rlabel metal3 s -960 373676 480 373916 4 la_data_out[99]
port 397 nsew signal tristate
rlabel metal3 s -960 339404 480 339644 4 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 469006 703520 469118 704960 6 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 455758 703520 455870 704960 6 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 555854 -960 555966 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 249494 -960 249606 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 56294 703520 56406 704960 6 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 562294 703520 562406 704960 6 la_oenb[104]
port 404 nsew signal input
rlabel metal3 s 583520 46732 584960 46972 6 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 465694 703520 465806 704960 6 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 142958 -960 143070 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal3 s -960 181916 480 182156 4 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 402766 -960 402878 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 538926 703520 539038 704960 6 la_oenb[10]
port 410 nsew signal input
rlabel metal3 s -960 614940 480 615180 4 la_oenb[110]
port 411 nsew signal input
rlabel metal3 s -960 693548 480 693788 4 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 432390 703520 432502 704960 6 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 219686 -960 219798 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal3 s 583520 558636 584960 558876 6 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 399270 -960 399382 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal3 s 583520 366604 584960 366844 6 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 329350 703520 329462 704960 6 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 319414 -960 319526 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 282798 -960 282910 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal3 s -960 344300 480 344540 4 la_oenb[120]
port 422 nsew signal input
rlabel metal3 s 583520 258348 584960 258588 6 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 82974 703520 83086 704960 6 la_oenb[122]
port 424 nsew signal input
rlabel metal3 s 583520 401148 584960 401388 6 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 149582 703520 149694 704960 6 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 196318 -960 196430 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 349222 703520 349334 704960 6 la_oenb[126]
port 428 nsew signal input
rlabel metal3 s -960 270588 480 270828 4 la_oenb[127]
port 429 nsew signal input
rlabel metal3 s 583520 214012 584960 214252 6 la_oenb[12]
port 430 nsew signal input
rlabel metal3 s 583520 332332 584960 332572 6 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 452630 -960 452742 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal3 s 583520 150092 584960 150332 6 la_oenb[15]
port 433 nsew signal input
rlabel metal3 s 583520 494716 584960 494956 6 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 345910 703520 346022 704960 6 la_oenb[17]
port 435 nsew signal input
rlabel metal3 s -960 186812 480 187052 4 la_oenb[18]
port 436 nsew signal input
rlabel metal3 s -960 88348 480 88588 4 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 156390 -960 156502 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal3 s 583520 86172 584960 86412 6 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 36606 -960 36718 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 163014 -960 163126 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal3 s 583520 66588 584960 66828 6 la_oenb[23]
port 442 nsew signal input
rlabel metal3 s 583520 686476 584960 686716 6 la_oenb[24]
port 443 nsew signal input
rlabel metal3 s 583520 278204 584960 278444 6 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 59790 -960 59902 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal3 s 583520 219180 584960 219420 6 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 379398 -960 379510 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 492374 703520 492486 704960 6 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 352718 -960 352830 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal3 s 583520 381564 584960 381804 6 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 558982 703520 559094 704960 6 la_oenb[31]
port 451 nsew signal input
rlabel metal3 s -960 280380 480 280620 4 la_oenb[32]
port 452 nsew signal input
rlabel metal3 s -960 600252 480 600492 4 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 565606 703520 565718 704960 6 la_oenb[34]
port 454 nsew signal input
rlabel metal3 s -960 117996 480 118236 4 la_oenb[35]
port 455 nsew signal input
rlabel metal3 s -960 368780 480 369020 4 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 582350 -960 582462 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal3 s -960 231148 480 231388 4 la_oenb[38]
port 458 nsew signal input
rlabel metal3 s -960 314652 480 314892 4 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 282614 703520 282726 704960 6 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 419326 -960 419438 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal3 s -960 477036 480 477276 4 la_oenb[41]
port 462 nsew signal input
rlabel metal3 s -960 408220 480 408460 4 la_oenb[42]
port 463 nsew signal input
rlabel metal3 s -960 403324 480 403564 4 la_oenb[43]
port 464 nsew signal input
rlabel metal3 s 583520 661996 584960 662236 6 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 502494 -960 502606 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal3 s -960 196604 480 196844 4 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 482622 -960 482734 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal3 s -960 191708 480 191948 4 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 96406 -960 96518 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 149766 -960 149878 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 519238 -960 519350 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal3 s 583520 184636 584960 184876 6 la_oenb[51]
port 473 nsew signal input
rlabel metal3 s 583520 592908 584960 593148 6 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 299358 703520 299470 704960 6 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 275990 703520 276102 704960 6 la_oenb[54]
port 476 nsew signal input
rlabel metal3 s -960 590188 480 590428 4 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 183070 -960 183182 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal3 s 583520 671788 584960 672028 6 la_oenb[57]
port 479 nsew signal input
rlabel metal3 s -960 358988 480 359228 4 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 159518 703520 159630 704960 6 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 116462 -960 116574 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal3 s 583520 578220 584960 578460 6 la_oenb[60]
port 483 nsew signal input
rlabel metal3 s -960 157164 480 157404 4 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 365966 703520 366078 704960 6 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 462382 703520 462494 704960 6 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 489062 703520 489174 704960 6 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 495686 703520 495798 704960 6 la_oenb[65]
port 488 nsew signal input
rlabel metal3 s -960 54076 480 54316 4 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 312606 703520 312718 704960 6 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 19862 -960 19974 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 6614 -960 6726 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal3 s -960 127788 480 128028 4 la_oenb[70]
port 494 nsew signal input
rlabel metal3 s 583520 95964 584960 96204 6 la_oenb[71]
port 495 nsew signal input
rlabel metal3 s -960 541228 480 541468 4 la_oenb[72]
port 496 nsew signal input
rlabel metal3 s -960 521372 480 521612 4 la_oenb[73]
port 497 nsew signal input
rlabel metal3 s -960 629628 480 629868 4 la_oenb[74]
port 498 nsew signal input
rlabel metal3 s -960 324716 480 324956 4 la_oenb[75]
port 499 nsew signal input
rlabel metal3 s -960 275484 480 275724 4 la_oenb[76]
port 500 nsew signal input
rlabel metal3 s -960 211292 480 211532 4 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 302670 703520 302782 704960 6 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 495870 -960 495982 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 236246 -960 236358 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal3 s -960 605148 480 605388 4 la_oenb[80]
port 505 nsew signal input
rlabel metal3 s 583520 489820 584960 490060 6 la_oenb[81]
port 506 nsew signal input
rlabel metal3 s 583520 652204 584960 652444 6 la_oenb[82]
port 507 nsew signal input
rlabel metal3 s -960 437868 480 438108 4 la_oenb[83]
port 508 nsew signal input
rlabel metal3 s -960 29324 480 29564 4 la_oenb[84]
port 509 nsew signal input
rlabel metal3 s 583520 32044 584960 32284 6 la_oenb[85]
port 510 nsew signal input
rlabel metal3 s 583520 612764 584960 613004 6 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 229438 703520 229550 704960 6 la_oenb[87]
port 512 nsew signal input
rlabel metal3 s 583520 499612 584960 499852 6 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 462566 -960 462678 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 362470 703520 362582 704960 6 la_oenb[8]
port 515 nsew signal input
rlabel metal3 s 583520 120716 584960 120956 6 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 189510 703520 189622 704960 6 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 559166 -960 559278 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal3 s -960 678860 480 679100 4 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 76534 -960 76646 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal3 s 583520 469964 584960 470204 6 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal3 s 583520 602972 584960 603212 6 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 153078 -960 153190 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 29614 703520 29726 704960 6 la_oenb[9]
port 526 nsew signal input
rlabel metal3 s -960 378844 480 379084 4 user_clock2
port 527 nsew signal input
rlabel metal3 s -960 172124 480 172364 4 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 9742 703520 9854 704960 6 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 62918 703520 63030 704960 6 user_irq[2]
port 530 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 wb_clk_i
port 531 nsew signal input
rlabel metal3 s -960 673964 480 674204 4 wb_rst_i
port 532 nsew signal input
rlabel metal3 s 583520 317372 584960 317612 6 wbs_ack_o
port 533 nsew signal tristate
rlabel metal2 s 266054 703520 266166 704960 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 142774 703520 142886 704960 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal3 s -960 575500 480 575740 4 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 53166 -960 53278 480 8 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal3 s -960 442764 480 443004 4 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal3 s 583520 642140 584960 642380 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal3 s 583520 588012 584960 588252 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal3 s 583520 524092 584960 524332 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal3 s 583520 273308 584960 273548 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 562478 -960 562590 480 8 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 272678 703520 272790 704960 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal3 s -960 255628 480 255868 4 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 329534 -960 329646 480 8 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 472502 -960 472614 480 8 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal3 s 583520 194428 584960 194668 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal3 s -960 669068 480 669308 4 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 316102 -960 316214 480 8 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 63102 -960 63214 480 8 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 109654 703520 109766 704960 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal3 s 583520 484652 584960 484892 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 515742 703520 515854 704960 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 222998 -960 223110 480 8 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 375902 703520 376014 704960 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal3 s 583520 347020 584960 347260 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 446006 -960 446118 480 8 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 369278 703520 369390 704960 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal3 s -960 132684 480 132924 4 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 179574 -960 179686 480 8 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 29798 -960 29910 480 8 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 572414 -960 572526 480 8 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal3 s 583520 209116 584960 209356 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 119590 703520 119702 704960 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 582166 703520 582278 704960 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal3 s -960 432972 480 433212 4 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal3 s -960 491996 480 492236 4 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal3 s -960 472140 480 472380 4 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 23174 -960 23286 480 8 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 123086 -960 123198 480 8 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal3 s 583520 406044 584960 406284 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal3 s -960 44012 480 44252 4 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 342598 703520 342710 704960 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 479126 703520 479238 704960 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal3 s -960 688652 480 688892 4 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 86470 -960 86582 480 8 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal3 s 583520 465068 584960 465308 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 498998 703520 499110 704960 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal3 s -960 319548 480 319788 4 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal3 s 583520 607868 584960 608108 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal3 s 583520 233868 584960 234108 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal3 s -960 19532 480 19772 4 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 439198 703520 439310 704960 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 112966 703520 113078 704960 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 176262 -960 176374 480 8 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal3 s 583520 455276 584960 455516 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 455942 -960 456054 480 8 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal3 s 583520 199324 584960 199564 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal3 s -960 299964 480 300204 4 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 575726 -960 575838 480 8 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 89782 -960 89894 480 8 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal3 s -960 4844 480 5084 4 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 429078 703520 429190 704960 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal3 s 583520 676684 584960 676924 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 579038 -960 579150 480 8 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 43230 -960 43342 480 8 wbs_dat_o[0]
port 599 nsew signal tristate
rlabel metal3 s 583520 410940 584960 411180 6 wbs_dat_o[10]
port 600 nsew signal tristate
rlabel metal2 s 13238 -960 13350 480 8 wbs_dat_o[11]
port 601 nsew signal tristate
rlabel metal3 s 583520 691372 584960 691612 6 wbs_dat_o[12]
port 602 nsew signal tristate
rlabel metal2 s 415830 703520 415942 704960 6 wbs_dat_o[13]
port 603 nsew signal tristate
rlabel metal3 s 583520 41836 584960 42076 6 wbs_dat_o[14]
port 604 nsew signal tristate
rlabel metal2 s 399086 703520 399198 704960 6 wbs_dat_o[15]
port 605 nsew signal tristate
rlabel metal2 s 369462 -960 369574 480 8 wbs_dat_o[16]
port 606 nsew signal tristate
rlabel metal3 s -960 14636 480 14876 4 wbs_dat_o[17]
port 607 nsew signal tristate
rlabel metal2 s 366150 -960 366262 480 8 wbs_dat_o[18]
port 608 nsew signal tristate
rlabel metal2 s -10 -960 102 480 8 wbs_dat_o[19]
port 609 nsew signal tristate
rlabel metal2 s 429262 -960 429374 480 8 wbs_dat_o[1]
port 610 nsew signal tristate
rlabel metal3 s -960 309756 480 309996 4 wbs_dat_o[20]
port 611 nsew signal tristate
rlabel metal3 s -960 624732 480 624972 4 wbs_dat_o[21]
port 612 nsew signal tristate
rlabel metal2 s 169454 703520 169566 704960 6 wbs_dat_o[22]
port 613 nsew signal tristate
rlabel metal3 s -960 201500 480 201740 4 wbs_dat_o[23]
port 614 nsew signal tristate
rlabel metal2 s 113150 -960 113262 480 8 wbs_dat_o[24]
port 615 nsew signal tristate
rlabel metal2 s 39918 -960 40030 480 8 wbs_dat_o[25]
port 616 nsew signal tristate
rlabel metal2 s 305982 703520 306094 704960 6 wbs_dat_o[26]
port 617 nsew signal tristate
rlabel metal2 s 186198 703520 186310 704960 6 wbs_dat_o[27]
port 618 nsew signal tristate
rlabel metal2 s 292918 -960 293030 480 8 wbs_dat_o[28]
port 619 nsew signal tristate
rlabel metal2 s 402582 703520 402694 704960 6 wbs_dat_o[29]
port 620 nsew signal tristate
rlabel metal3 s 583520 154988 584960 155228 6 wbs_dat_o[2]
port 621 nsew signal tristate
rlabel metal3 s -960 481932 480 482172 4 wbs_dat_o[30]
port 622 nsew signal tristate
rlabel metal3 s 583520 543948 584960 544188 6 wbs_dat_o[31]
port 623 nsew signal tristate
rlabel metal2 s 119774 -960 119886 480 8 wbs_dat_o[3]
port 624 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 wbs_dat_o[4]
port 625 nsew signal tristate
rlabel metal2 s 322726 -960 322838 480 8 wbs_dat_o[5]
port 626 nsew signal tristate
rlabel metal3 s 583520 509404 584960 509644 6 wbs_dat_o[6]
port 627 nsew signal tristate
rlabel metal2 s 326038 -960 326150 480 8 wbs_dat_o[7]
port 628 nsew signal tristate
rlabel metal2 s 392462 703520 392574 704960 6 wbs_dat_o[8]
port 629 nsew signal tristate
rlabel metal2 s 389150 703520 389262 704960 6 wbs_dat_o[9]
port 630 nsew signal tristate
rlabel metal2 s 6430 703520 6542 704960 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 102846 703520 102958 704960 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 386022 -960 386134 480 8 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal3 s -960 167228 480 167468 4 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal3 s -960 644316 480 644556 4 wbs_stb_i
port 635 nsew signal input
rlabel metal3 s 583520 307580 584960 307820 6 wbs_we_i
port 636 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
