VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 3100.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.790 -4.800 2256.350 2.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 -4.800 136.670 2.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1229.180 2504.800 1230.380 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 738.220 2.400 739.420 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.630 3097.600 947.190 3104.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1945.900 2504.800 1947.100 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.110 3097.600 826.670 3104.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2953.660 2504.800 2954.860 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1140.780 2.400 1141.980 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.990 3097.600 1023.550 3104.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 -4.800 212.110 2.400 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.750 3097.600 750.310 3104.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 3097.600 871.750 3104.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 312.540 2.400 313.740 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 849.740 2.400 850.940 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2236.940 2504.800 2238.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 3097.600 250.750 3104.800 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.350 3097.600 1628.910 3104.800 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.750 3097.600 796.310 3104.800 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 133.020 2.400 134.220 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.870 3097.600 1220.430 3104.800 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2775.500 2.400 2776.700 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.430 -4.800 983.990 2.400 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 984.380 2.400 985.580 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.790 3097.600 1750.350 3104.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.550 3097.600 1523.110 3104.800 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.390 -4.800 696.950 2.400 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1967.660 2504.800 1968.860 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1162.540 2.400 1163.740 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.270 -4.800 2135.830 2.400 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1185.660 2.400 1186.860 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.790 3097.600 2371.350 3104.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 154.780 2504.800 155.980 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1721.500 2504.800 1722.700 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1879.260 2.400 1880.460 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.670 3097.600 1280.230 3104.800 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2193.420 2.400 2194.620 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 938.140 2504.800 939.340 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 871.500 2504.800 872.700 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.910 3097.600 1553.470 3104.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.990 3097.600 977.550 3104.800 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.150 -4.800 1711.710 2.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.510 3097.600 569.070 3104.800 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 959.900 2504.800 961.100 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.070 -4.800 1574.630 2.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 3097.600 175.310 3104.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 3097.600 220.390 3104.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1029.260 2.400 1030.460 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.350 -4.800 1559.910 2.400 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.230 3097.600 583.790 3104.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.510 3097.600 1765.070 3104.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 603.580 2.400 604.780 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1117.660 2504.800 1118.860 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 3065.180 2504.800 3066.380 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2640.860 2.400 2642.060 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.350 3097.600 432.910 3104.800 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 43.260 2.400 44.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.270 3097.600 1583.830 3104.800 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2213.820 2504.800 2215.020 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2639.500 2504.800 2640.700 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.910 -4.800 1438.470 2.400 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2976.780 2.400 2977.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.790 3097.600 462.350 3104.800 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 3097.600 265.470 3104.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.870 3097.600 599.430 3104.800 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1834.380 2.400 1835.580 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.430 -4.800 1029.990 2.400 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2484.460 2.400 2485.660 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.670 3097.600 1947.230 3104.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.590 -4.800 1166.150 2.400 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 916.380 2.400 917.580 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 3097.600 1840.510 3104.800 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.870 3097.600 2416.430 3104.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2394.700 2.400 2395.900 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.990 3097.600 402.550 3104.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 3097.600 144.950 3104.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 3097.600 2355.710 3104.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2863.900 2504.800 2865.100 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1095.900 2.400 1097.100 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 2.400 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2348.460 2504.800 2349.660 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 512.460 2504.800 513.660 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1922.780 2504.800 1923.980 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2751.020 2504.800 2752.220 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2371.580 2504.800 2372.780 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 -4.800 272.830 2.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.950 -4.800 1771.510 2.400 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 3097.600 114.590 3104.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.070 -4.800 2195.630 2.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 109.900 2504.800 111.100 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2304.940 2.400 2306.140 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 3097.600 629.790 3104.800 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.510 -4.800 2317.070 2.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1609.980 2504.800 1611.180 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.590 -4.800 545.150 2.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2401.150 3097.600 2401.710 3104.800 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.750 -4.800 727.310 2.400 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2706.140 2504.800 2707.340 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2281.820 2504.800 2283.020 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.590 3097.600 2477.150 3104.800 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2012.540 2504.800 2013.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.590 3097.600 614.150 3104.800 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2074.550 -4.800 2075.110 2.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1656.220 2.400 1657.420 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 65.020 2504.800 66.220 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1833.020 2504.800 1834.220 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 3097.600 1340.950 3104.800 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 783.100 2.400 784.300 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.150 3097.600 1113.710 3104.800 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 3097.600 129.310 3104.800 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1094.540 2504.800 1095.740 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.390 3097.600 2007.950 3104.800 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1453.580 2504.800 1454.780 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 691.980 2504.800 693.180 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.510 3097.600 1190.070 3104.800 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.150 3097.600 538.710 3104.800 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2819.020 2504.800 2820.220 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2551.100 2.400 2552.300 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1856.140 2504.800 1857.340 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 86.780 2504.800 87.980 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.470 3097.600 1432.030 3104.800 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 625.340 2504.800 626.540 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.230 3097.600 1825.790 3104.800 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2617.740 2.400 2618.940 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.390 -4.800 75.950 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1877.900 2504.800 1879.100 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2662.620 2.400 2663.820 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 266.300 2504.800 267.500 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.950 3097.600 1886.510 3104.800 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.230 -4.800 560.790 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 -4.800 1014.350 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.430 3097.600 1098.990 3104.800 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.830 3097.600 2037.390 3104.800 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1766.380 2504.800 1767.580 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2439.580 2.400 2440.780 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.150 3097.600 1734.710 3104.800 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.070 -4.800 2241.630 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 3097.600 281.110 3104.800 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2346.870 -4.800 2347.430 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.630 3097.600 372.190 3104.800 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 871.500 2.400 872.700 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.230 -4.800 1756.790 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1812.620 2.400 1813.820 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1521.580 2.400 1522.780 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.190 -4.800 2044.750 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2168.940 2504.800 2170.140 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 536.940 2.400 538.140 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1162.540 2504.800 1163.740 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1386.940 2.400 1388.140 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2572.860 2504.800 2574.060 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.030 3097.600 1931.590 3104.800 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.950 -4.800 575.510 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 3097.600 205.670 3104.800 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 111.260 2.400 112.460 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.990 -4.800 1529.550 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1520.220 2504.800 1521.420 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 400.940 2504.800 402.140 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2238.300 2.400 2239.500 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2438.220 2504.800 2439.420 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 245.900 2.400 247.100 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1744.620 2504.800 1745.820 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.430 -4.800 1650.990 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.670 -4.800 1832.230 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.710 -4.800 2165.270 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 3097.600 1007.910 3104.800 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.790 -4.800 1681.350 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.590 3097.600 1235.150 3104.800 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2820.380 2.400 2821.580 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.750 3097.600 1992.310 3104.800 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2430.590 3097.600 2431.150 3104.800 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1207.420 2504.800 1208.620 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 -4.800 45.590 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1744.620 2.400 1745.820 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.150 -4.800 469.710 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1274.060 2504.800 1275.260 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2326.700 2504.800 2327.900 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.910 3097.600 932.470 3104.800 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 580.460 2.400 581.660 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1857.500 2.400 1858.700 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.630 -4.800 1545.190 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 3097.600 1811.070 3104.800 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.510 -4.800 454.070 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.190 -4.800 802.750 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 66.380 2.400 67.580 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 3097.600 190.030 3104.800 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2385.510 3097.600 2386.070 3104.800 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 377.820 2504.800 379.020 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.990 -4.800 287.550 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 -4.800 15.230 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.870 -4.800 1726.430 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.550 3097.600 2098.110 3104.800 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.830 -4.800 2014.390 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1431.820 2.400 1433.020 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 3097.600 341.830 3104.800 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.870 -4.800 484.430 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 557.340 2504.800 558.540 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2908.780 2504.800 2909.980 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.190 -4.800 1998.750 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 3097.600 53.870 3104.800 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.790 3097.600 1129.350 3104.800 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 827.980 2.400 829.180 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2192.060 2504.800 2193.260 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1072.780 2504.800 1073.980 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 580.460 2504.800 581.660 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 356.060 2504.800 357.260 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.030 3097.600 735.590 3104.800 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.230 -4.800 1135.790 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.990 -4.800 908.550 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1901.020 2504.800 1902.220 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2415.100 2504.800 2416.300 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 668.860 2504.800 670.060 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 781.740 2504.800 782.940 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.390 -4.800 1892.950 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 803.500 2504.800 804.700 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1498.460 2.400 1499.660 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.190 3097.600 2113.750 3104.800 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 21.500 2.400 22.700 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.790 3097.600 1083.350 3104.800 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2124.060 2504.800 2125.260 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1701.100 2.400 1702.300 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2058.780 2.400 2059.980 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.270 3097.600 962.830 3104.800 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.670 3097.600 705.230 3104.800 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.910 3097.600 1507.470 3104.800 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 3097.600 236.030 3104.800 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.590 -4.800 2362.150 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.910 -4.800 817.470 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.630 -4.800 924.190 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 20.140 2504.800 21.340 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1207.420 2.400 1208.620 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2953.660 2.400 2954.860 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1318.940 2504.800 1320.140 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2283.180 2.400 2284.380 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.430 -4.800 408.990 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2125.420 2.400 2126.620 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.790 3097.600 2325.350 3104.800 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2931.900 2.400 2933.100 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 289.420 2.400 290.620 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 983.020 2504.800 984.220 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1565.100 2504.800 1566.300 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3097.600 689.590 3104.800 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.270 -4.800 1514.830 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2685.740 2.400 2686.940 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.750 3097.600 1371.310 3104.800 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.630 3097.600 1568.190 3104.800 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.350 -4.800 363.910 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 3097.600 1870.870 3104.800 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.710 3097.600 2280.270 3104.800 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 267.660 2.400 268.860 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 3097.600 1144.070 3104.800 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2684.380 2504.800 2685.580 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 490.700 2504.800 491.900 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 804.860 2.400 806.060 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.630 -4.800 878.190 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1230.540 2.400 1231.740 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.390 -4.800 1317.950 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2391.950 -4.800 2392.510 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.870 3097.600 553.430 3104.800 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 3097.600 2310.630 3104.800 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2707.500 2.400 2708.700 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1119.020 2.400 1120.220 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.910 -4.800 2105.470 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.110 -4.800 1332.670 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2035.660 2.400 2036.860 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2729.260 2504.800 2730.460 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1250.940 2504.800 1252.140 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1320.300 2.400 1321.500 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1408.700 2504.800 1409.900 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2271.430 -4.800 2271.990 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.990 3097.600 356.550 3104.800 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 311.180 2504.800 312.380 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2170.300 2.400 2171.500 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.630 3097.600 326.190 3104.800 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2997.180 2504.800 2998.380 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 693.340 2.400 694.540 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.070 3097.600 1689.630 3104.800 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1004.780 2504.800 1005.980 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.790 -4.800 1060.350 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.830 3097.600 1462.390 3104.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 670.220 2.400 671.420 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1295.820 2504.800 1297.020 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 -4.800 348.270 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 3097.600 23.510 3104.800 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 221.420 2504.800 222.620 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.510 -4.800 1075.070 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1006.140 2.400 1007.340 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 3097.600 659.230 3104.800 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 3097.600 1492.750 3104.800 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.430 -4.800 2225.990 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 3097.600 2219.550 3104.800 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2529.340 2.400 2530.540 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1611.340 2.400 1612.540 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.110 3097.600 2022.670 3104.800 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 647.100 2504.800 648.300 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.430 3097.600 1052.990 3104.800 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2148.540 2.400 2149.740 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.750 -4.800 1302.310 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.910 3097.600 886.470 3104.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.470 3097.600 811.030 3104.800 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.390 -4.800 1938.950 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.230 -4.800 2377.790 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.950 3097.600 2461.510 3104.800 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.630 3097.600 993.190 3104.800 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 402.300 2.400 403.500 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.470 -4.800 167.030 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1588.220 2.400 1589.420 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1924.140 2.400 1925.340 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.110 -4.800 711.670 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2574.220 2.400 2575.420 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1430.460 2504.800 1431.660 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2080.540 2.400 2081.740 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1340.700 2504.800 1341.900 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 177.900 2.400 179.100 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.670 -4.800 1211.230 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.430 3097.600 2340.990 3104.800 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.390 3097.600 1961.950 3104.800 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.310 3097.600 1295.870 3104.800 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.350 -4.800 317.910 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.950 -4.800 1817.510 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2887.020 2.400 2888.220 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1541.980 2504.800 1543.180 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 467.580 2504.800 468.780 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 176.540 2504.800 177.740 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.870 -4.800 1105.430 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.790 -4.800 1635.350 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.270 -4.800 847.830 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.070 3097.600 2264.630 3104.800 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.670 -4.800 1257.230 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.070 3097.600 1068.630 3104.800 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 3097.600 68.590 3104.800 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.030 -4.800 620.590 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.670 3097.600 1326.230 3104.800 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.870 -4.800 1151.430 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 43.260 2504.800 44.460 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.350 -4.800 2180.910 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 445.820 2504.800 447.020 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 289.420 2504.800 290.620 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.910 -4.800 863.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 3097.600 8.790 3104.800 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 424.060 2.400 425.260 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.310 3097.600 674.870 3104.800 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.670 -4.800 1878.230 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 3097.600 508.350 3104.800 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 625.340 2.400 626.540 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1475.340 2504.800 1476.540 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.190 3097.600 1446.750 3104.800 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.390 3097.600 1386.950 3104.800 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.110 3097.600 1401.670 3104.800 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.510 -4.800 1742.070 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 3097.600 2144.110 3104.800 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.270 3097.600 916.830 3104.800 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.150 3097.600 1159.710 3104.800 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.310 -4.800 1801.870 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.350 3097.600 386.910 3104.800 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1275.420 2.400 1276.620 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.830 3097.600 2083.390 3104.800 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.150 -4.800 2332.710 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.150 -4.800 1044.710 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.310 -4.800 1226.870 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 3042.060 2504.800 3043.260 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2842.140 2.400 2843.340 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.910 3097.600 2128.470 3104.800 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.670 -4.800 590.230 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1676.620 2504.800 1677.820 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.310 3097.600 1249.870 3104.800 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.230 3097.600 2446.790 3104.800 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1631.740 2504.800 1632.940 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.790 3097.600 1704.350 3104.800 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.030 3097.600 1977.590 3104.800 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.350 -4.800 938.910 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2303.580 2504.800 2304.780 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.510 -4.800 1696.070 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1767.740 2.400 1768.940 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.790 -4.800 439.350 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.270 3097.600 1537.830 3104.800 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.750 -4.800 1348.310 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.950 -4.800 1196.510 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2930.540 2504.800 2931.740 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1049.660 2504.800 1050.860 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1633.100 2.400 1634.300 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1654.860 2504.800 1656.060 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.910 -4.800 1484.470 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.550 -4.800 833.110 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2461.340 2.400 2462.540 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2527.980 2504.800 2529.180 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1969.020 2.400 1970.220 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2326.700 2.400 2327.900 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.030 -4.800 1908.590 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 602.220 2504.800 603.420 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2057.420 2504.800 2058.620 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 558.700 2.400 559.900 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 468.940 2.400 470.140 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.030 -4.800 1241.590 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.030 -4.800 666.590 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 334.300 2504.800 335.500 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 -4.800 151.390 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.750 -4.800 681.310 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 244.540 2504.800 245.740 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2885.660 2504.800 2886.860 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1139.420 2504.800 1140.620 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.910 -4.800 242.470 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1051.020 2.400 1052.220 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.270 3097.600 2204.830 3104.800 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.630 -4.800 1499.190 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1586.860 2504.800 1588.060 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.310 3097.600 2491.870 3104.800 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2233.710 3097.600 2234.270 3104.800 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 156.140 2.400 157.340 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1566.460 2.400 1567.660 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 3097.600 841.390 3104.800 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.830 -4.800 772.390 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.070 3097.600 447.630 3104.800 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 826.620 2504.800 827.820 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1699.740 2504.800 1700.940 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 447.180 2.400 448.380 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2483.100 2504.800 2484.300 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2260.060 2.400 2261.260 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.430 3097.600 2294.990 3104.800 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.780 2.400 2909.980 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.990 -4.800 2150.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.270 3097.600 295.830 3104.800 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2865.260 2.400 2866.460 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2468.310 -4.800 2468.870 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.150 -4.800 423.710 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.670 -4.800 636.230 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.710 -4.800 2211.270 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 758.620 2504.800 759.820 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2504.860 2504.800 2506.060 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2349.820 2.400 2351.020 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.950 3097.600 1265.510 3104.800 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.550 3097.600 902.110 3104.800 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1677.980 2.400 1679.180 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2840.780 2504.800 2841.980 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2506.220 2.400 2507.420 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.390 3097.600 765.950 3104.800 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 492.060 2.400 493.260 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2459.980 2504.800 2461.180 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.870 3097.600 1795.430 3104.800 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 3097.600 39.150 3104.800 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.470 3097.600 2053.030 3104.800 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.910 3097.600 2174.470 3104.800 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.630 3097.600 2189.190 3104.800 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.190 -4.800 1377.750 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.750 3097.600 1417.310 3104.800 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 -4.800 90.670 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 -4.800 29.950 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.910 -4.800 2059.470 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1410.060 2.400 1411.260 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 422.700 2504.800 423.900 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1789.500 2.400 1790.700 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2371.580 2.400 2372.780 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 3097.600 98.950 3104.800 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1476.700 2.400 1477.900 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1252.300 2.400 1253.500 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 961.260 2.400 962.460 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 3097.600 1356.590 3104.800 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.070 -4.800 999.630 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2752.380 2.400 2753.580 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2080.540 2504.800 2081.740 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2795.900 2504.800 2797.100 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1992.140 2.400 1993.340 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2416.460 2.400 2417.660 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 131.660 2504.800 132.860 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2617.740 2504.800 2618.940 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.710 3097.600 1038.270 3104.800 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2147.180 2504.800 2148.380 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.470 -4.800 1984.030 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1722.860 2.400 1724.060 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 535.580 2504.800 536.780 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.550 3097.600 856.110 3104.800 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.590 -4.800 2408.150 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3066.540 2.400 3067.740 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.990 -4.800 333.550 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1297.180 2.400 1298.380 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2594.620 2504.800 2595.820 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.390 -4.800 650.950 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.110 3097.600 159.670 3104.800 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.630 3097.600 1614.190 3104.800 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 513.820 2.400 515.020 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 3097.600 84.230 3104.800 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.910 3097.600 311.470 3104.800 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 736.860 2504.800 738.060 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3021.660 2.400 3022.860 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 939.500 2.400 940.700 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 3097.600 1174.430 3104.800 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.950 3097.600 644.510 3104.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2595.980 2.400 2597.180 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.270 -4.800 226.830 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2013.900 2.400 2015.100 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2774.140 2504.800 2775.340 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2549.740 2504.800 2550.940 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 222.780 2.400 223.980 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1184.300 2504.800 1185.500 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.310 -4.800 2422.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.230 3097.600 1204.790 3104.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.310 3097.600 1916.870 3104.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.190 -4.800 1423.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.550 -4.800 2029.110 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 848.380 2504.800 849.580 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2998.540 2.400 2999.740 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.470 -4.800 1363.030 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.150 3097.600 492.710 3104.800 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2102.300 2504.800 2103.500 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2249.350 3097.600 2249.910 3104.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.710 -4.800 969.270 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.070 3097.600 1643.630 3104.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1498.460 2504.800 1499.660 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.750 -4.800 1923.310 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.990 3097.600 1598.550 3104.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.310 -4.800 1847.870 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.550 -4.800 787.110 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 -4.800 121.030 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 916.380 2504.800 917.580 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 3097.600 523.070 3104.800 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 3086.940 2504.800 3088.140 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1947.260 2.400 1948.460 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2215.180 2.400 2216.380 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 334.300 2.400 335.500 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.750 -4.800 106.310 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.870 -4.800 530.430 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1789.500 2504.800 1790.700 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.830 -4.800 1393.390 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.550 3097.600 1477.110 3104.800 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.190 3097.600 2067.750 3104.800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3043.420 2.400 3044.620 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.070 -4.800 378.630 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2035.660 2504.800 2036.860 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.270 3097.600 2158.830 3104.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1453.580 2.400 1454.780 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2662.620 2504.800 2663.820 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1027.900 2504.800 1029.100 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 88.140 2.400 89.340 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.670 3097.600 1901.230 3104.800 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.430 3097.600 477.990 3104.800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.110 -4.800 757.670 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1990.780 2504.800 1991.980 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.830 -4.800 1968.390 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 893.260 2504.800 894.460 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1342.060 2.400 1343.260 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.030 -4.800 2483.590 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.310 -4.800 1180.870 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1363.820 2504.800 1365.020 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.590 3097.600 1856.150 3104.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2975.420 2504.800 2976.620 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.670 -4.800 2499.230 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.910 -4.800 196.470 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1811.260 2504.800 1812.460 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 -4.800 60.310 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 3020.300 2504.800 3021.500 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.150 3097.600 1780.710 3104.800 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 199.660 2504.800 200.860 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 379.180 2.400 380.380 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 648.460 2.400 649.660 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 759.980 2.400 761.180 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.710 -4.800 1590.270 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 -4.800 0.510 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.030 -4.800 1862.590 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1365.180 2.400 1366.380 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2730.620 2.400 2731.820 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.390 3097.600 719.950 3104.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 894.620 2.400 895.820 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.510 -4.800 500.070 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 -4.800 181.750 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.030 3097.600 1310.590 3104.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.110 3097.600 780.670 3104.800 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.390 -4.800 1271.950 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.430 3097.600 1719.990 3104.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 713.740 2504.800 714.940 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2103.660 2.400 2104.860 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2393.340 2504.800 2394.540 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.230 -4.800 514.790 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.270 -4.800 893.830 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 201.020 2.400 202.220 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 2258.700 2504.800 2259.900 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.550 -4.800 1408.110 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.430 3097.600 1673.990 3104.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.710 3097.600 1659.270 3104.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3088.300 2.400 3089.500 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.710 3097.600 417.270 3104.800 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.150 -4.800 1665.710 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 715.100 2.400 716.300 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2797.260 2.400 2798.460 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2497.600 1385.580 2504.800 1386.780 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 15.180 15.045 2491.215 3076.405 ;
      LAYER met1 ;
        RECT 0.070 13.980 2499.110 3087.840 ;
      LAYER met2 ;
        RECT 0.100 3097.320 7.950 3097.810 ;
        RECT 9.070 3097.320 22.670 3097.810 ;
        RECT 23.790 3097.320 38.310 3097.810 ;
        RECT 39.430 3097.320 53.030 3097.810 ;
        RECT 54.150 3097.320 67.750 3097.810 ;
        RECT 68.870 3097.320 83.390 3097.810 ;
        RECT 84.510 3097.320 98.110 3097.810 ;
        RECT 99.230 3097.320 113.750 3097.810 ;
        RECT 114.870 3097.320 128.470 3097.810 ;
        RECT 129.590 3097.320 144.110 3097.810 ;
        RECT 145.230 3097.320 158.830 3097.810 ;
        RECT 159.950 3097.320 174.470 3097.810 ;
        RECT 175.590 3097.320 189.190 3097.810 ;
        RECT 190.310 3097.320 204.830 3097.810 ;
        RECT 205.950 3097.320 219.550 3097.810 ;
        RECT 220.670 3097.320 235.190 3097.810 ;
        RECT 236.310 3097.320 249.910 3097.810 ;
        RECT 251.030 3097.320 264.630 3097.810 ;
        RECT 265.750 3097.320 280.270 3097.810 ;
        RECT 281.390 3097.320 294.990 3097.810 ;
        RECT 296.110 3097.320 310.630 3097.810 ;
        RECT 311.750 3097.320 325.350 3097.810 ;
        RECT 326.470 3097.320 340.990 3097.810 ;
        RECT 342.110 3097.320 355.710 3097.810 ;
        RECT 356.830 3097.320 371.350 3097.810 ;
        RECT 372.470 3097.320 386.070 3097.810 ;
        RECT 387.190 3097.320 401.710 3097.810 ;
        RECT 402.830 3097.320 416.430 3097.810 ;
        RECT 417.550 3097.320 432.070 3097.810 ;
        RECT 433.190 3097.320 446.790 3097.810 ;
        RECT 447.910 3097.320 461.510 3097.810 ;
        RECT 462.630 3097.320 477.150 3097.810 ;
        RECT 478.270 3097.320 491.870 3097.810 ;
        RECT 492.990 3097.320 507.510 3097.810 ;
        RECT 508.630 3097.320 522.230 3097.810 ;
        RECT 523.350 3097.320 537.870 3097.810 ;
        RECT 538.990 3097.320 552.590 3097.810 ;
        RECT 553.710 3097.320 568.230 3097.810 ;
        RECT 569.350 3097.320 582.950 3097.810 ;
        RECT 584.070 3097.320 598.590 3097.810 ;
        RECT 599.710 3097.320 613.310 3097.810 ;
        RECT 614.430 3097.320 628.950 3097.810 ;
        RECT 630.070 3097.320 643.670 3097.810 ;
        RECT 644.790 3097.320 658.390 3097.810 ;
        RECT 659.510 3097.320 674.030 3097.810 ;
        RECT 675.150 3097.320 688.750 3097.810 ;
        RECT 689.870 3097.320 704.390 3097.810 ;
        RECT 705.510 3097.320 719.110 3097.810 ;
        RECT 720.230 3097.320 734.750 3097.810 ;
        RECT 735.870 3097.320 749.470 3097.810 ;
        RECT 750.590 3097.320 765.110 3097.810 ;
        RECT 766.230 3097.320 779.830 3097.810 ;
        RECT 780.950 3097.320 795.470 3097.810 ;
        RECT 796.590 3097.320 810.190 3097.810 ;
        RECT 811.310 3097.320 825.830 3097.810 ;
        RECT 826.950 3097.320 840.550 3097.810 ;
        RECT 841.670 3097.320 855.270 3097.810 ;
        RECT 856.390 3097.320 870.910 3097.810 ;
        RECT 872.030 3097.320 885.630 3097.810 ;
        RECT 886.750 3097.320 901.270 3097.810 ;
        RECT 902.390 3097.320 915.990 3097.810 ;
        RECT 917.110 3097.320 931.630 3097.810 ;
        RECT 932.750 3097.320 946.350 3097.810 ;
        RECT 947.470 3097.320 961.990 3097.810 ;
        RECT 963.110 3097.320 976.710 3097.810 ;
        RECT 977.830 3097.320 992.350 3097.810 ;
        RECT 993.470 3097.320 1007.070 3097.810 ;
        RECT 1008.190 3097.320 1022.710 3097.810 ;
        RECT 1023.830 3097.320 1037.430 3097.810 ;
        RECT 1038.550 3097.320 1052.150 3097.810 ;
        RECT 1053.270 3097.320 1067.790 3097.810 ;
        RECT 1068.910 3097.320 1082.510 3097.810 ;
        RECT 1083.630 3097.320 1098.150 3097.810 ;
        RECT 1099.270 3097.320 1112.870 3097.810 ;
        RECT 1113.990 3097.320 1128.510 3097.810 ;
        RECT 1129.630 3097.320 1143.230 3097.810 ;
        RECT 1144.350 3097.320 1158.870 3097.810 ;
        RECT 1159.990 3097.320 1173.590 3097.810 ;
        RECT 1174.710 3097.320 1189.230 3097.810 ;
        RECT 1190.350 3097.320 1203.950 3097.810 ;
        RECT 1205.070 3097.320 1219.590 3097.810 ;
        RECT 1220.710 3097.320 1234.310 3097.810 ;
        RECT 1235.430 3097.320 1249.030 3097.810 ;
        RECT 1250.150 3097.320 1264.670 3097.810 ;
        RECT 1265.790 3097.320 1279.390 3097.810 ;
        RECT 1280.510 3097.320 1295.030 3097.810 ;
        RECT 1296.150 3097.320 1309.750 3097.810 ;
        RECT 1310.870 3097.320 1325.390 3097.810 ;
        RECT 1326.510 3097.320 1340.110 3097.810 ;
        RECT 1341.230 3097.320 1355.750 3097.810 ;
        RECT 1356.870 3097.320 1370.470 3097.810 ;
        RECT 1371.590 3097.320 1386.110 3097.810 ;
        RECT 1387.230 3097.320 1400.830 3097.810 ;
        RECT 1401.950 3097.320 1416.470 3097.810 ;
        RECT 1417.590 3097.320 1431.190 3097.810 ;
        RECT 1432.310 3097.320 1445.910 3097.810 ;
        RECT 1447.030 3097.320 1461.550 3097.810 ;
        RECT 1462.670 3097.320 1476.270 3097.810 ;
        RECT 1477.390 3097.320 1491.910 3097.810 ;
        RECT 1493.030 3097.320 1506.630 3097.810 ;
        RECT 1507.750 3097.320 1522.270 3097.810 ;
        RECT 1523.390 3097.320 1536.990 3097.810 ;
        RECT 1538.110 3097.320 1552.630 3097.810 ;
        RECT 1553.750 3097.320 1567.350 3097.810 ;
        RECT 1568.470 3097.320 1582.990 3097.810 ;
        RECT 1584.110 3097.320 1597.710 3097.810 ;
        RECT 1598.830 3097.320 1613.350 3097.810 ;
        RECT 1614.470 3097.320 1628.070 3097.810 ;
        RECT 1629.190 3097.320 1642.790 3097.810 ;
        RECT 1643.910 3097.320 1658.430 3097.810 ;
        RECT 1659.550 3097.320 1673.150 3097.810 ;
        RECT 1674.270 3097.320 1688.790 3097.810 ;
        RECT 1689.910 3097.320 1703.510 3097.810 ;
        RECT 1704.630 3097.320 1719.150 3097.810 ;
        RECT 1720.270 3097.320 1733.870 3097.810 ;
        RECT 1734.990 3097.320 1749.510 3097.810 ;
        RECT 1750.630 3097.320 1764.230 3097.810 ;
        RECT 1765.350 3097.320 1779.870 3097.810 ;
        RECT 1780.990 3097.320 1794.590 3097.810 ;
        RECT 1795.710 3097.320 1810.230 3097.810 ;
        RECT 1811.350 3097.320 1824.950 3097.810 ;
        RECT 1826.070 3097.320 1839.670 3097.810 ;
        RECT 1840.790 3097.320 1855.310 3097.810 ;
        RECT 1856.430 3097.320 1870.030 3097.810 ;
        RECT 1871.150 3097.320 1885.670 3097.810 ;
        RECT 1886.790 3097.320 1900.390 3097.810 ;
        RECT 1901.510 3097.320 1916.030 3097.810 ;
        RECT 1917.150 3097.320 1930.750 3097.810 ;
        RECT 1931.870 3097.320 1946.390 3097.810 ;
        RECT 1947.510 3097.320 1961.110 3097.810 ;
        RECT 1962.230 3097.320 1976.750 3097.810 ;
        RECT 1977.870 3097.320 1991.470 3097.810 ;
        RECT 1992.590 3097.320 2007.110 3097.810 ;
        RECT 2008.230 3097.320 2021.830 3097.810 ;
        RECT 2022.950 3097.320 2036.550 3097.810 ;
        RECT 2037.670 3097.320 2052.190 3097.810 ;
        RECT 2053.310 3097.320 2066.910 3097.810 ;
        RECT 2068.030 3097.320 2082.550 3097.810 ;
        RECT 2083.670 3097.320 2097.270 3097.810 ;
        RECT 2098.390 3097.320 2112.910 3097.810 ;
        RECT 2114.030 3097.320 2127.630 3097.810 ;
        RECT 2128.750 3097.320 2143.270 3097.810 ;
        RECT 2144.390 3097.320 2157.990 3097.810 ;
        RECT 2159.110 3097.320 2173.630 3097.810 ;
        RECT 2174.750 3097.320 2188.350 3097.810 ;
        RECT 2189.470 3097.320 2203.990 3097.810 ;
        RECT 2205.110 3097.320 2218.710 3097.810 ;
        RECT 2219.830 3097.320 2233.430 3097.810 ;
        RECT 2234.550 3097.320 2249.070 3097.810 ;
        RECT 2250.190 3097.320 2263.790 3097.810 ;
        RECT 2264.910 3097.320 2279.430 3097.810 ;
        RECT 2280.550 3097.320 2294.150 3097.810 ;
        RECT 2295.270 3097.320 2309.790 3097.810 ;
        RECT 2310.910 3097.320 2324.510 3097.810 ;
        RECT 2325.630 3097.320 2340.150 3097.810 ;
        RECT 2341.270 3097.320 2354.870 3097.810 ;
        RECT 2355.990 3097.320 2370.510 3097.810 ;
        RECT 2371.630 3097.320 2385.230 3097.810 ;
        RECT 2386.350 3097.320 2400.870 3097.810 ;
        RECT 2401.990 3097.320 2415.590 3097.810 ;
        RECT 2416.710 3097.320 2430.310 3097.810 ;
        RECT 2431.430 3097.320 2445.950 3097.810 ;
        RECT 2447.070 3097.320 2460.670 3097.810 ;
        RECT 2461.790 3097.320 2476.310 3097.810 ;
        RECT 2477.430 3097.320 2491.030 3097.810 ;
        RECT 2492.150 3097.320 2499.080 3097.810 ;
        RECT 0.100 2.680 2499.080 3097.320 ;
        RECT 0.790 2.310 14.390 2.680 ;
        RECT 15.510 2.310 29.110 2.680 ;
        RECT 30.230 2.310 44.750 2.680 ;
        RECT 45.870 2.310 59.470 2.680 ;
        RECT 60.590 2.310 75.110 2.680 ;
        RECT 76.230 2.310 89.830 2.680 ;
        RECT 90.950 2.310 105.470 2.680 ;
        RECT 106.590 2.310 120.190 2.680 ;
        RECT 121.310 2.310 135.830 2.680 ;
        RECT 136.950 2.310 150.550 2.680 ;
        RECT 151.670 2.310 166.190 2.680 ;
        RECT 167.310 2.310 180.910 2.680 ;
        RECT 182.030 2.310 195.630 2.680 ;
        RECT 196.750 2.310 211.270 2.680 ;
        RECT 212.390 2.310 225.990 2.680 ;
        RECT 227.110 2.310 241.630 2.680 ;
        RECT 242.750 2.310 256.350 2.680 ;
        RECT 257.470 2.310 271.990 2.680 ;
        RECT 273.110 2.310 286.710 2.680 ;
        RECT 287.830 2.310 302.350 2.680 ;
        RECT 303.470 2.310 317.070 2.680 ;
        RECT 318.190 2.310 332.710 2.680 ;
        RECT 333.830 2.310 347.430 2.680 ;
        RECT 348.550 2.310 363.070 2.680 ;
        RECT 364.190 2.310 377.790 2.680 ;
        RECT 378.910 2.310 392.510 2.680 ;
        RECT 393.630 2.310 408.150 2.680 ;
        RECT 409.270 2.310 422.870 2.680 ;
        RECT 423.990 2.310 438.510 2.680 ;
        RECT 439.630 2.310 453.230 2.680 ;
        RECT 454.350 2.310 468.870 2.680 ;
        RECT 469.990 2.310 483.590 2.680 ;
        RECT 484.710 2.310 499.230 2.680 ;
        RECT 500.350 2.310 513.950 2.680 ;
        RECT 515.070 2.310 529.590 2.680 ;
        RECT 530.710 2.310 544.310 2.680 ;
        RECT 545.430 2.310 559.950 2.680 ;
        RECT 561.070 2.310 574.670 2.680 ;
        RECT 575.790 2.310 589.390 2.680 ;
        RECT 590.510 2.310 605.030 2.680 ;
        RECT 606.150 2.310 619.750 2.680 ;
        RECT 620.870 2.310 635.390 2.680 ;
        RECT 636.510 2.310 650.110 2.680 ;
        RECT 651.230 2.310 665.750 2.680 ;
        RECT 666.870 2.310 680.470 2.680 ;
        RECT 681.590 2.310 696.110 2.680 ;
        RECT 697.230 2.310 710.830 2.680 ;
        RECT 711.950 2.310 726.470 2.680 ;
        RECT 727.590 2.310 741.190 2.680 ;
        RECT 742.310 2.310 756.830 2.680 ;
        RECT 757.950 2.310 771.550 2.680 ;
        RECT 772.670 2.310 786.270 2.680 ;
        RECT 787.390 2.310 801.910 2.680 ;
        RECT 803.030 2.310 816.630 2.680 ;
        RECT 817.750 2.310 832.270 2.680 ;
        RECT 833.390 2.310 846.990 2.680 ;
        RECT 848.110 2.310 862.630 2.680 ;
        RECT 863.750 2.310 877.350 2.680 ;
        RECT 878.470 2.310 892.990 2.680 ;
        RECT 894.110 2.310 907.710 2.680 ;
        RECT 908.830 2.310 923.350 2.680 ;
        RECT 924.470 2.310 938.070 2.680 ;
        RECT 939.190 2.310 953.710 2.680 ;
        RECT 954.830 2.310 968.430 2.680 ;
        RECT 969.550 2.310 983.150 2.680 ;
        RECT 984.270 2.310 998.790 2.680 ;
        RECT 999.910 2.310 1013.510 2.680 ;
        RECT 1014.630 2.310 1029.150 2.680 ;
        RECT 1030.270 2.310 1043.870 2.680 ;
        RECT 1044.990 2.310 1059.510 2.680 ;
        RECT 1060.630 2.310 1074.230 2.680 ;
        RECT 1075.350 2.310 1089.870 2.680 ;
        RECT 1090.990 2.310 1104.590 2.680 ;
        RECT 1105.710 2.310 1120.230 2.680 ;
        RECT 1121.350 2.310 1134.950 2.680 ;
        RECT 1136.070 2.310 1150.590 2.680 ;
        RECT 1151.710 2.310 1165.310 2.680 ;
        RECT 1166.430 2.310 1180.030 2.680 ;
        RECT 1181.150 2.310 1195.670 2.680 ;
        RECT 1196.790 2.310 1210.390 2.680 ;
        RECT 1211.510 2.310 1226.030 2.680 ;
        RECT 1227.150 2.310 1240.750 2.680 ;
        RECT 1241.870 2.310 1256.390 2.680 ;
        RECT 1257.510 2.310 1271.110 2.680 ;
        RECT 1272.230 2.310 1286.750 2.680 ;
        RECT 1287.870 2.310 1301.470 2.680 ;
        RECT 1302.590 2.310 1317.110 2.680 ;
        RECT 1318.230 2.310 1331.830 2.680 ;
        RECT 1332.950 2.310 1347.470 2.680 ;
        RECT 1348.590 2.310 1362.190 2.680 ;
        RECT 1363.310 2.310 1376.910 2.680 ;
        RECT 1378.030 2.310 1392.550 2.680 ;
        RECT 1393.670 2.310 1407.270 2.680 ;
        RECT 1408.390 2.310 1422.910 2.680 ;
        RECT 1424.030 2.310 1437.630 2.680 ;
        RECT 1438.750 2.310 1453.270 2.680 ;
        RECT 1454.390 2.310 1467.990 2.680 ;
        RECT 1469.110 2.310 1483.630 2.680 ;
        RECT 1484.750 2.310 1498.350 2.680 ;
        RECT 1499.470 2.310 1513.990 2.680 ;
        RECT 1515.110 2.310 1528.710 2.680 ;
        RECT 1529.830 2.310 1544.350 2.680 ;
        RECT 1545.470 2.310 1559.070 2.680 ;
        RECT 1560.190 2.310 1573.790 2.680 ;
        RECT 1574.910 2.310 1589.430 2.680 ;
        RECT 1590.550 2.310 1604.150 2.680 ;
        RECT 1605.270 2.310 1619.790 2.680 ;
        RECT 1620.910 2.310 1634.510 2.680 ;
        RECT 1635.630 2.310 1650.150 2.680 ;
        RECT 1651.270 2.310 1664.870 2.680 ;
        RECT 1665.990 2.310 1680.510 2.680 ;
        RECT 1681.630 2.310 1695.230 2.680 ;
        RECT 1696.350 2.310 1710.870 2.680 ;
        RECT 1711.990 2.310 1725.590 2.680 ;
        RECT 1726.710 2.310 1741.230 2.680 ;
        RECT 1742.350 2.310 1755.950 2.680 ;
        RECT 1757.070 2.310 1770.670 2.680 ;
        RECT 1771.790 2.310 1786.310 2.680 ;
        RECT 1787.430 2.310 1801.030 2.680 ;
        RECT 1802.150 2.310 1816.670 2.680 ;
        RECT 1817.790 2.310 1831.390 2.680 ;
        RECT 1832.510 2.310 1847.030 2.680 ;
        RECT 1848.150 2.310 1861.750 2.680 ;
        RECT 1862.870 2.310 1877.390 2.680 ;
        RECT 1878.510 2.310 1892.110 2.680 ;
        RECT 1893.230 2.310 1907.750 2.680 ;
        RECT 1908.870 2.310 1922.470 2.680 ;
        RECT 1923.590 2.310 1938.110 2.680 ;
        RECT 1939.230 2.310 1952.830 2.680 ;
        RECT 1953.950 2.310 1967.550 2.680 ;
        RECT 1968.670 2.310 1983.190 2.680 ;
        RECT 1984.310 2.310 1997.910 2.680 ;
        RECT 1999.030 2.310 2013.550 2.680 ;
        RECT 2014.670 2.310 2028.270 2.680 ;
        RECT 2029.390 2.310 2043.910 2.680 ;
        RECT 2045.030 2.310 2058.630 2.680 ;
        RECT 2059.750 2.310 2074.270 2.680 ;
        RECT 2075.390 2.310 2088.990 2.680 ;
        RECT 2090.110 2.310 2104.630 2.680 ;
        RECT 2105.750 2.310 2119.350 2.680 ;
        RECT 2120.470 2.310 2134.990 2.680 ;
        RECT 2136.110 2.310 2149.710 2.680 ;
        RECT 2150.830 2.310 2164.430 2.680 ;
        RECT 2165.550 2.310 2180.070 2.680 ;
        RECT 2181.190 2.310 2194.790 2.680 ;
        RECT 2195.910 2.310 2210.430 2.680 ;
        RECT 2211.550 2.310 2225.150 2.680 ;
        RECT 2226.270 2.310 2240.790 2.680 ;
        RECT 2241.910 2.310 2255.510 2.680 ;
        RECT 2256.630 2.310 2271.150 2.680 ;
        RECT 2272.270 2.310 2285.870 2.680 ;
        RECT 2286.990 2.310 2301.510 2.680 ;
        RECT 2302.630 2.310 2316.230 2.680 ;
        RECT 2317.350 2.310 2331.870 2.680 ;
        RECT 2332.990 2.310 2346.590 2.680 ;
        RECT 2347.710 2.310 2361.310 2.680 ;
        RECT 2362.430 2.310 2376.950 2.680 ;
        RECT 2378.070 2.310 2391.670 2.680 ;
        RECT 2392.790 2.310 2407.310 2.680 ;
        RECT 2408.430 2.310 2422.030 2.680 ;
        RECT 2423.150 2.310 2437.670 2.680 ;
        RECT 2438.790 2.310 2452.390 2.680 ;
        RECT 2453.510 2.310 2468.030 2.680 ;
        RECT 2469.150 2.310 2482.750 2.680 ;
        RECT 2483.870 2.310 2498.390 2.680 ;
      LAYER met3 ;
        RECT 2.800 3088.540 2497.600 3089.065 ;
        RECT 2.800 3087.900 2497.200 3088.540 ;
        RECT 2.400 3086.540 2497.200 3087.900 ;
        RECT 2.400 3068.140 2497.600 3086.540 ;
        RECT 2.800 3066.780 2497.600 3068.140 ;
        RECT 2.800 3066.140 2497.200 3066.780 ;
        RECT 2.400 3064.780 2497.200 3066.140 ;
        RECT 2.400 3045.020 2497.600 3064.780 ;
        RECT 2.800 3043.660 2497.600 3045.020 ;
        RECT 2.800 3043.020 2497.200 3043.660 ;
        RECT 2.400 3041.660 2497.200 3043.020 ;
        RECT 2.400 3023.260 2497.600 3041.660 ;
        RECT 2.800 3021.900 2497.600 3023.260 ;
        RECT 2.800 3021.260 2497.200 3021.900 ;
        RECT 2.400 3019.900 2497.200 3021.260 ;
        RECT 2.400 3000.140 2497.600 3019.900 ;
        RECT 2.800 2998.780 2497.600 3000.140 ;
        RECT 2.800 2998.140 2497.200 2998.780 ;
        RECT 2.400 2996.780 2497.200 2998.140 ;
        RECT 2.400 2978.380 2497.600 2996.780 ;
        RECT 2.800 2977.020 2497.600 2978.380 ;
        RECT 2.800 2976.380 2497.200 2977.020 ;
        RECT 2.400 2975.020 2497.200 2976.380 ;
        RECT 2.400 2955.260 2497.600 2975.020 ;
        RECT 2.800 2953.260 2497.200 2955.260 ;
        RECT 2.400 2933.500 2497.600 2953.260 ;
        RECT 2.800 2932.140 2497.600 2933.500 ;
        RECT 2.800 2931.500 2497.200 2932.140 ;
        RECT 2.400 2930.140 2497.200 2931.500 ;
        RECT 2.400 2910.380 2497.600 2930.140 ;
        RECT 2.800 2908.380 2497.200 2910.380 ;
        RECT 2.400 2888.620 2497.600 2908.380 ;
        RECT 2.800 2887.260 2497.600 2888.620 ;
        RECT 2.800 2886.620 2497.200 2887.260 ;
        RECT 2.400 2885.260 2497.200 2886.620 ;
        RECT 2.400 2866.860 2497.600 2885.260 ;
        RECT 2.800 2865.500 2497.600 2866.860 ;
        RECT 2.800 2864.860 2497.200 2865.500 ;
        RECT 2.400 2863.500 2497.200 2864.860 ;
        RECT 2.400 2843.740 2497.600 2863.500 ;
        RECT 2.800 2842.380 2497.600 2843.740 ;
        RECT 2.800 2841.740 2497.200 2842.380 ;
        RECT 2.400 2840.380 2497.200 2841.740 ;
        RECT 2.400 2821.980 2497.600 2840.380 ;
        RECT 2.800 2820.620 2497.600 2821.980 ;
        RECT 2.800 2819.980 2497.200 2820.620 ;
        RECT 2.400 2818.620 2497.200 2819.980 ;
        RECT 2.400 2798.860 2497.600 2818.620 ;
        RECT 2.800 2797.500 2497.600 2798.860 ;
        RECT 2.800 2796.860 2497.200 2797.500 ;
        RECT 2.400 2795.500 2497.200 2796.860 ;
        RECT 2.400 2777.100 2497.600 2795.500 ;
        RECT 2.800 2775.740 2497.600 2777.100 ;
        RECT 2.800 2775.100 2497.200 2775.740 ;
        RECT 2.400 2773.740 2497.200 2775.100 ;
        RECT 2.400 2753.980 2497.600 2773.740 ;
        RECT 2.800 2752.620 2497.600 2753.980 ;
        RECT 2.800 2751.980 2497.200 2752.620 ;
        RECT 2.400 2750.620 2497.200 2751.980 ;
        RECT 2.400 2732.220 2497.600 2750.620 ;
        RECT 2.800 2730.860 2497.600 2732.220 ;
        RECT 2.800 2730.220 2497.200 2730.860 ;
        RECT 2.400 2728.860 2497.200 2730.220 ;
        RECT 2.400 2709.100 2497.600 2728.860 ;
        RECT 2.800 2707.740 2497.600 2709.100 ;
        RECT 2.800 2707.100 2497.200 2707.740 ;
        RECT 2.400 2705.740 2497.200 2707.100 ;
        RECT 2.400 2687.340 2497.600 2705.740 ;
        RECT 2.800 2685.980 2497.600 2687.340 ;
        RECT 2.800 2685.340 2497.200 2685.980 ;
        RECT 2.400 2683.980 2497.200 2685.340 ;
        RECT 2.400 2664.220 2497.600 2683.980 ;
        RECT 2.800 2662.220 2497.200 2664.220 ;
        RECT 2.400 2642.460 2497.600 2662.220 ;
        RECT 2.800 2641.100 2497.600 2642.460 ;
        RECT 2.800 2640.460 2497.200 2641.100 ;
        RECT 2.400 2639.100 2497.200 2640.460 ;
        RECT 2.400 2619.340 2497.600 2639.100 ;
        RECT 2.800 2617.340 2497.200 2619.340 ;
        RECT 2.400 2597.580 2497.600 2617.340 ;
        RECT 2.800 2596.220 2497.600 2597.580 ;
        RECT 2.800 2595.580 2497.200 2596.220 ;
        RECT 2.400 2594.220 2497.200 2595.580 ;
        RECT 2.400 2575.820 2497.600 2594.220 ;
        RECT 2.800 2574.460 2497.600 2575.820 ;
        RECT 2.800 2573.820 2497.200 2574.460 ;
        RECT 2.400 2572.460 2497.200 2573.820 ;
        RECT 2.400 2552.700 2497.600 2572.460 ;
        RECT 2.800 2551.340 2497.600 2552.700 ;
        RECT 2.800 2550.700 2497.200 2551.340 ;
        RECT 2.400 2549.340 2497.200 2550.700 ;
        RECT 2.400 2530.940 2497.600 2549.340 ;
        RECT 2.800 2529.580 2497.600 2530.940 ;
        RECT 2.800 2528.940 2497.200 2529.580 ;
        RECT 2.400 2527.580 2497.200 2528.940 ;
        RECT 2.400 2507.820 2497.600 2527.580 ;
        RECT 2.800 2506.460 2497.600 2507.820 ;
        RECT 2.800 2505.820 2497.200 2506.460 ;
        RECT 2.400 2504.460 2497.200 2505.820 ;
        RECT 2.400 2486.060 2497.600 2504.460 ;
        RECT 2.800 2484.700 2497.600 2486.060 ;
        RECT 2.800 2484.060 2497.200 2484.700 ;
        RECT 2.400 2482.700 2497.200 2484.060 ;
        RECT 2.400 2462.940 2497.600 2482.700 ;
        RECT 2.800 2461.580 2497.600 2462.940 ;
        RECT 2.800 2460.940 2497.200 2461.580 ;
        RECT 2.400 2459.580 2497.200 2460.940 ;
        RECT 2.400 2441.180 2497.600 2459.580 ;
        RECT 2.800 2439.820 2497.600 2441.180 ;
        RECT 2.800 2439.180 2497.200 2439.820 ;
        RECT 2.400 2437.820 2497.200 2439.180 ;
        RECT 2.400 2418.060 2497.600 2437.820 ;
        RECT 2.800 2416.700 2497.600 2418.060 ;
        RECT 2.800 2416.060 2497.200 2416.700 ;
        RECT 2.400 2414.700 2497.200 2416.060 ;
        RECT 2.400 2396.300 2497.600 2414.700 ;
        RECT 2.800 2394.940 2497.600 2396.300 ;
        RECT 2.800 2394.300 2497.200 2394.940 ;
        RECT 2.400 2392.940 2497.200 2394.300 ;
        RECT 2.400 2373.180 2497.600 2392.940 ;
        RECT 2.800 2371.180 2497.200 2373.180 ;
        RECT 2.400 2351.420 2497.600 2371.180 ;
        RECT 2.800 2350.060 2497.600 2351.420 ;
        RECT 2.800 2349.420 2497.200 2350.060 ;
        RECT 2.400 2348.060 2497.200 2349.420 ;
        RECT 2.400 2328.300 2497.600 2348.060 ;
        RECT 2.800 2326.300 2497.200 2328.300 ;
        RECT 2.400 2306.540 2497.600 2326.300 ;
        RECT 2.800 2305.180 2497.600 2306.540 ;
        RECT 2.800 2304.540 2497.200 2305.180 ;
        RECT 2.400 2303.180 2497.200 2304.540 ;
        RECT 2.400 2284.780 2497.600 2303.180 ;
        RECT 2.800 2283.420 2497.600 2284.780 ;
        RECT 2.800 2282.780 2497.200 2283.420 ;
        RECT 2.400 2281.420 2497.200 2282.780 ;
        RECT 2.400 2261.660 2497.600 2281.420 ;
        RECT 2.800 2260.300 2497.600 2261.660 ;
        RECT 2.800 2259.660 2497.200 2260.300 ;
        RECT 2.400 2258.300 2497.200 2259.660 ;
        RECT 2.400 2239.900 2497.600 2258.300 ;
        RECT 2.800 2238.540 2497.600 2239.900 ;
        RECT 2.800 2237.900 2497.200 2238.540 ;
        RECT 2.400 2236.540 2497.200 2237.900 ;
        RECT 2.400 2216.780 2497.600 2236.540 ;
        RECT 2.800 2215.420 2497.600 2216.780 ;
        RECT 2.800 2214.780 2497.200 2215.420 ;
        RECT 2.400 2213.420 2497.200 2214.780 ;
        RECT 2.400 2195.020 2497.600 2213.420 ;
        RECT 2.800 2193.660 2497.600 2195.020 ;
        RECT 2.800 2193.020 2497.200 2193.660 ;
        RECT 2.400 2191.660 2497.200 2193.020 ;
        RECT 2.400 2171.900 2497.600 2191.660 ;
        RECT 2.800 2170.540 2497.600 2171.900 ;
        RECT 2.800 2169.900 2497.200 2170.540 ;
        RECT 2.400 2168.540 2497.200 2169.900 ;
        RECT 2.400 2150.140 2497.600 2168.540 ;
        RECT 2.800 2148.780 2497.600 2150.140 ;
        RECT 2.800 2148.140 2497.200 2148.780 ;
        RECT 2.400 2146.780 2497.200 2148.140 ;
        RECT 2.400 2127.020 2497.600 2146.780 ;
        RECT 2.800 2125.660 2497.600 2127.020 ;
        RECT 2.800 2125.020 2497.200 2125.660 ;
        RECT 2.400 2123.660 2497.200 2125.020 ;
        RECT 2.400 2105.260 2497.600 2123.660 ;
        RECT 2.800 2103.900 2497.600 2105.260 ;
        RECT 2.800 2103.260 2497.200 2103.900 ;
        RECT 2.400 2101.900 2497.200 2103.260 ;
        RECT 2.400 2082.140 2497.600 2101.900 ;
        RECT 2.800 2080.140 2497.200 2082.140 ;
        RECT 2.400 2060.380 2497.600 2080.140 ;
        RECT 2.800 2059.020 2497.600 2060.380 ;
        RECT 2.800 2058.380 2497.200 2059.020 ;
        RECT 2.400 2057.020 2497.200 2058.380 ;
        RECT 2.400 2037.260 2497.600 2057.020 ;
        RECT 2.800 2035.260 2497.200 2037.260 ;
        RECT 2.400 2015.500 2497.600 2035.260 ;
        RECT 2.800 2014.140 2497.600 2015.500 ;
        RECT 2.800 2013.500 2497.200 2014.140 ;
        RECT 2.400 2012.140 2497.200 2013.500 ;
        RECT 2.400 1993.740 2497.600 2012.140 ;
        RECT 2.800 1992.380 2497.600 1993.740 ;
        RECT 2.800 1991.740 2497.200 1992.380 ;
        RECT 2.400 1990.380 2497.200 1991.740 ;
        RECT 2.400 1970.620 2497.600 1990.380 ;
        RECT 2.800 1969.260 2497.600 1970.620 ;
        RECT 2.800 1968.620 2497.200 1969.260 ;
        RECT 2.400 1967.260 2497.200 1968.620 ;
        RECT 2.400 1948.860 2497.600 1967.260 ;
        RECT 2.800 1947.500 2497.600 1948.860 ;
        RECT 2.800 1946.860 2497.200 1947.500 ;
        RECT 2.400 1945.500 2497.200 1946.860 ;
        RECT 2.400 1925.740 2497.600 1945.500 ;
        RECT 2.800 1924.380 2497.600 1925.740 ;
        RECT 2.800 1923.740 2497.200 1924.380 ;
        RECT 2.400 1922.380 2497.200 1923.740 ;
        RECT 2.400 1903.980 2497.600 1922.380 ;
        RECT 2.800 1902.620 2497.600 1903.980 ;
        RECT 2.800 1901.980 2497.200 1902.620 ;
        RECT 2.400 1900.620 2497.200 1901.980 ;
        RECT 2.400 1880.860 2497.600 1900.620 ;
        RECT 2.800 1879.500 2497.600 1880.860 ;
        RECT 2.800 1878.860 2497.200 1879.500 ;
        RECT 2.400 1877.500 2497.200 1878.860 ;
        RECT 2.400 1859.100 2497.600 1877.500 ;
        RECT 2.800 1857.740 2497.600 1859.100 ;
        RECT 2.800 1857.100 2497.200 1857.740 ;
        RECT 2.400 1855.740 2497.200 1857.100 ;
        RECT 2.400 1835.980 2497.600 1855.740 ;
        RECT 2.800 1834.620 2497.600 1835.980 ;
        RECT 2.800 1833.980 2497.200 1834.620 ;
        RECT 2.400 1832.620 2497.200 1833.980 ;
        RECT 2.400 1814.220 2497.600 1832.620 ;
        RECT 2.800 1812.860 2497.600 1814.220 ;
        RECT 2.800 1812.220 2497.200 1812.860 ;
        RECT 2.400 1810.860 2497.200 1812.220 ;
        RECT 2.400 1791.100 2497.600 1810.860 ;
        RECT 2.800 1789.100 2497.200 1791.100 ;
        RECT 2.400 1769.340 2497.600 1789.100 ;
        RECT 2.800 1767.980 2497.600 1769.340 ;
        RECT 2.800 1767.340 2497.200 1767.980 ;
        RECT 2.400 1765.980 2497.200 1767.340 ;
        RECT 2.400 1746.220 2497.600 1765.980 ;
        RECT 2.800 1744.220 2497.200 1746.220 ;
        RECT 2.400 1724.460 2497.600 1744.220 ;
        RECT 2.800 1723.100 2497.600 1724.460 ;
        RECT 2.800 1722.460 2497.200 1723.100 ;
        RECT 2.400 1721.100 2497.200 1722.460 ;
        RECT 2.400 1702.700 2497.600 1721.100 ;
        RECT 2.800 1701.340 2497.600 1702.700 ;
        RECT 2.800 1700.700 2497.200 1701.340 ;
        RECT 2.400 1699.340 2497.200 1700.700 ;
        RECT 2.400 1679.580 2497.600 1699.340 ;
        RECT 2.800 1678.220 2497.600 1679.580 ;
        RECT 2.800 1677.580 2497.200 1678.220 ;
        RECT 2.400 1676.220 2497.200 1677.580 ;
        RECT 2.400 1657.820 2497.600 1676.220 ;
        RECT 2.800 1656.460 2497.600 1657.820 ;
        RECT 2.800 1655.820 2497.200 1656.460 ;
        RECT 2.400 1654.460 2497.200 1655.820 ;
        RECT 2.400 1634.700 2497.600 1654.460 ;
        RECT 2.800 1633.340 2497.600 1634.700 ;
        RECT 2.800 1632.700 2497.200 1633.340 ;
        RECT 2.400 1631.340 2497.200 1632.700 ;
        RECT 2.400 1612.940 2497.600 1631.340 ;
        RECT 2.800 1611.580 2497.600 1612.940 ;
        RECT 2.800 1610.940 2497.200 1611.580 ;
        RECT 2.400 1609.580 2497.200 1610.940 ;
        RECT 2.400 1589.820 2497.600 1609.580 ;
        RECT 2.800 1588.460 2497.600 1589.820 ;
        RECT 2.800 1587.820 2497.200 1588.460 ;
        RECT 2.400 1586.460 2497.200 1587.820 ;
        RECT 2.400 1568.060 2497.600 1586.460 ;
        RECT 2.800 1566.700 2497.600 1568.060 ;
        RECT 2.800 1566.060 2497.200 1566.700 ;
        RECT 2.400 1564.700 2497.200 1566.060 ;
        RECT 2.400 1544.940 2497.600 1564.700 ;
        RECT 2.800 1543.580 2497.600 1544.940 ;
        RECT 2.800 1542.940 2497.200 1543.580 ;
        RECT 2.400 1541.580 2497.200 1542.940 ;
        RECT 2.400 1523.180 2497.600 1541.580 ;
        RECT 2.800 1521.820 2497.600 1523.180 ;
        RECT 2.800 1521.180 2497.200 1521.820 ;
        RECT 2.400 1519.820 2497.200 1521.180 ;
        RECT 2.400 1500.060 2497.600 1519.820 ;
        RECT 2.800 1498.060 2497.200 1500.060 ;
        RECT 2.400 1478.300 2497.600 1498.060 ;
        RECT 2.800 1476.940 2497.600 1478.300 ;
        RECT 2.800 1476.300 2497.200 1476.940 ;
        RECT 2.400 1474.940 2497.200 1476.300 ;
        RECT 2.400 1455.180 2497.600 1474.940 ;
        RECT 2.800 1453.180 2497.200 1455.180 ;
        RECT 2.400 1433.420 2497.600 1453.180 ;
        RECT 2.800 1432.060 2497.600 1433.420 ;
        RECT 2.800 1431.420 2497.200 1432.060 ;
        RECT 2.400 1430.060 2497.200 1431.420 ;
        RECT 2.400 1411.660 2497.600 1430.060 ;
        RECT 2.800 1410.300 2497.600 1411.660 ;
        RECT 2.800 1409.660 2497.200 1410.300 ;
        RECT 2.400 1408.300 2497.200 1409.660 ;
        RECT 2.400 1388.540 2497.600 1408.300 ;
        RECT 2.800 1387.180 2497.600 1388.540 ;
        RECT 2.800 1386.540 2497.200 1387.180 ;
        RECT 2.400 1385.180 2497.200 1386.540 ;
        RECT 2.400 1366.780 2497.600 1385.180 ;
        RECT 2.800 1365.420 2497.600 1366.780 ;
        RECT 2.800 1364.780 2497.200 1365.420 ;
        RECT 2.400 1363.420 2497.200 1364.780 ;
        RECT 2.400 1343.660 2497.600 1363.420 ;
        RECT 2.800 1342.300 2497.600 1343.660 ;
        RECT 2.800 1341.660 2497.200 1342.300 ;
        RECT 2.400 1340.300 2497.200 1341.660 ;
        RECT 2.400 1321.900 2497.600 1340.300 ;
        RECT 2.800 1320.540 2497.600 1321.900 ;
        RECT 2.800 1319.900 2497.200 1320.540 ;
        RECT 2.400 1318.540 2497.200 1319.900 ;
        RECT 2.400 1298.780 2497.600 1318.540 ;
        RECT 2.800 1297.420 2497.600 1298.780 ;
        RECT 2.800 1296.780 2497.200 1297.420 ;
        RECT 2.400 1295.420 2497.200 1296.780 ;
        RECT 2.400 1277.020 2497.600 1295.420 ;
        RECT 2.800 1275.660 2497.600 1277.020 ;
        RECT 2.800 1275.020 2497.200 1275.660 ;
        RECT 2.400 1273.660 2497.200 1275.020 ;
        RECT 2.400 1253.900 2497.600 1273.660 ;
        RECT 2.800 1252.540 2497.600 1253.900 ;
        RECT 2.800 1251.900 2497.200 1252.540 ;
        RECT 2.400 1250.540 2497.200 1251.900 ;
        RECT 2.400 1232.140 2497.600 1250.540 ;
        RECT 2.800 1230.780 2497.600 1232.140 ;
        RECT 2.800 1230.140 2497.200 1230.780 ;
        RECT 2.400 1228.780 2497.200 1230.140 ;
        RECT 2.400 1209.020 2497.600 1228.780 ;
        RECT 2.800 1207.020 2497.200 1209.020 ;
        RECT 2.400 1187.260 2497.600 1207.020 ;
        RECT 2.800 1185.900 2497.600 1187.260 ;
        RECT 2.800 1185.260 2497.200 1185.900 ;
        RECT 2.400 1183.900 2497.200 1185.260 ;
        RECT 2.400 1164.140 2497.600 1183.900 ;
        RECT 2.800 1162.140 2497.200 1164.140 ;
        RECT 2.400 1142.380 2497.600 1162.140 ;
        RECT 2.800 1141.020 2497.600 1142.380 ;
        RECT 2.800 1140.380 2497.200 1141.020 ;
        RECT 2.400 1139.020 2497.200 1140.380 ;
        RECT 2.400 1120.620 2497.600 1139.020 ;
        RECT 2.800 1119.260 2497.600 1120.620 ;
        RECT 2.800 1118.620 2497.200 1119.260 ;
        RECT 2.400 1117.260 2497.200 1118.620 ;
        RECT 2.400 1097.500 2497.600 1117.260 ;
        RECT 2.800 1096.140 2497.600 1097.500 ;
        RECT 2.800 1095.500 2497.200 1096.140 ;
        RECT 2.400 1094.140 2497.200 1095.500 ;
        RECT 2.400 1075.740 2497.600 1094.140 ;
        RECT 2.800 1074.380 2497.600 1075.740 ;
        RECT 2.800 1073.740 2497.200 1074.380 ;
        RECT 2.400 1072.380 2497.200 1073.740 ;
        RECT 2.400 1052.620 2497.600 1072.380 ;
        RECT 2.800 1051.260 2497.600 1052.620 ;
        RECT 2.800 1050.620 2497.200 1051.260 ;
        RECT 2.400 1049.260 2497.200 1050.620 ;
        RECT 2.400 1030.860 2497.600 1049.260 ;
        RECT 2.800 1029.500 2497.600 1030.860 ;
        RECT 2.800 1028.860 2497.200 1029.500 ;
        RECT 2.400 1027.500 2497.200 1028.860 ;
        RECT 2.400 1007.740 2497.600 1027.500 ;
        RECT 2.800 1006.380 2497.600 1007.740 ;
        RECT 2.800 1005.740 2497.200 1006.380 ;
        RECT 2.400 1004.380 2497.200 1005.740 ;
        RECT 2.400 985.980 2497.600 1004.380 ;
        RECT 2.800 984.620 2497.600 985.980 ;
        RECT 2.800 983.980 2497.200 984.620 ;
        RECT 2.400 982.620 2497.200 983.980 ;
        RECT 2.400 962.860 2497.600 982.620 ;
        RECT 2.800 961.500 2497.600 962.860 ;
        RECT 2.800 960.860 2497.200 961.500 ;
        RECT 2.400 959.500 2497.200 960.860 ;
        RECT 2.400 941.100 2497.600 959.500 ;
        RECT 2.800 939.740 2497.600 941.100 ;
        RECT 2.800 939.100 2497.200 939.740 ;
        RECT 2.400 937.740 2497.200 939.100 ;
        RECT 2.400 917.980 2497.600 937.740 ;
        RECT 2.800 915.980 2497.200 917.980 ;
        RECT 2.400 896.220 2497.600 915.980 ;
        RECT 2.800 894.860 2497.600 896.220 ;
        RECT 2.800 894.220 2497.200 894.860 ;
        RECT 2.400 892.860 2497.200 894.220 ;
        RECT 2.400 873.100 2497.600 892.860 ;
        RECT 2.800 871.100 2497.200 873.100 ;
        RECT 2.400 851.340 2497.600 871.100 ;
        RECT 2.800 849.980 2497.600 851.340 ;
        RECT 2.800 849.340 2497.200 849.980 ;
        RECT 2.400 847.980 2497.200 849.340 ;
        RECT 2.400 829.580 2497.600 847.980 ;
        RECT 2.800 828.220 2497.600 829.580 ;
        RECT 2.800 827.580 2497.200 828.220 ;
        RECT 2.400 826.220 2497.200 827.580 ;
        RECT 2.400 806.460 2497.600 826.220 ;
        RECT 2.800 805.100 2497.600 806.460 ;
        RECT 2.800 804.460 2497.200 805.100 ;
        RECT 2.400 803.100 2497.200 804.460 ;
        RECT 2.400 784.700 2497.600 803.100 ;
        RECT 2.800 783.340 2497.600 784.700 ;
        RECT 2.800 782.700 2497.200 783.340 ;
        RECT 2.400 781.340 2497.200 782.700 ;
        RECT 2.400 761.580 2497.600 781.340 ;
        RECT 2.800 760.220 2497.600 761.580 ;
        RECT 2.800 759.580 2497.200 760.220 ;
        RECT 2.400 758.220 2497.200 759.580 ;
        RECT 2.400 739.820 2497.600 758.220 ;
        RECT 2.800 738.460 2497.600 739.820 ;
        RECT 2.800 737.820 2497.200 738.460 ;
        RECT 2.400 736.460 2497.200 737.820 ;
        RECT 2.400 716.700 2497.600 736.460 ;
        RECT 2.800 715.340 2497.600 716.700 ;
        RECT 2.800 714.700 2497.200 715.340 ;
        RECT 2.400 713.340 2497.200 714.700 ;
        RECT 2.400 694.940 2497.600 713.340 ;
        RECT 2.800 693.580 2497.600 694.940 ;
        RECT 2.800 692.940 2497.200 693.580 ;
        RECT 2.400 691.580 2497.200 692.940 ;
        RECT 2.400 671.820 2497.600 691.580 ;
        RECT 2.800 670.460 2497.600 671.820 ;
        RECT 2.800 669.820 2497.200 670.460 ;
        RECT 2.400 668.460 2497.200 669.820 ;
        RECT 2.400 650.060 2497.600 668.460 ;
        RECT 2.800 648.700 2497.600 650.060 ;
        RECT 2.800 648.060 2497.200 648.700 ;
        RECT 2.400 646.700 2497.200 648.060 ;
        RECT 2.400 626.940 2497.600 646.700 ;
        RECT 2.800 624.940 2497.200 626.940 ;
        RECT 2.400 605.180 2497.600 624.940 ;
        RECT 2.800 603.820 2497.600 605.180 ;
        RECT 2.800 603.180 2497.200 603.820 ;
        RECT 2.400 601.820 2497.200 603.180 ;
        RECT 2.400 582.060 2497.600 601.820 ;
        RECT 2.800 580.060 2497.200 582.060 ;
        RECT 2.400 560.300 2497.600 580.060 ;
        RECT 2.800 558.940 2497.600 560.300 ;
        RECT 2.800 558.300 2497.200 558.940 ;
        RECT 2.400 556.940 2497.200 558.300 ;
        RECT 2.400 538.540 2497.600 556.940 ;
        RECT 2.800 537.180 2497.600 538.540 ;
        RECT 2.800 536.540 2497.200 537.180 ;
        RECT 2.400 535.180 2497.200 536.540 ;
        RECT 2.400 515.420 2497.600 535.180 ;
        RECT 2.800 514.060 2497.600 515.420 ;
        RECT 2.800 513.420 2497.200 514.060 ;
        RECT 2.400 512.060 2497.200 513.420 ;
        RECT 2.400 493.660 2497.600 512.060 ;
        RECT 2.800 492.300 2497.600 493.660 ;
        RECT 2.800 491.660 2497.200 492.300 ;
        RECT 2.400 490.300 2497.200 491.660 ;
        RECT 2.400 470.540 2497.600 490.300 ;
        RECT 2.800 469.180 2497.600 470.540 ;
        RECT 2.800 468.540 2497.200 469.180 ;
        RECT 2.400 467.180 2497.200 468.540 ;
        RECT 2.400 448.780 2497.600 467.180 ;
        RECT 2.800 447.420 2497.600 448.780 ;
        RECT 2.800 446.780 2497.200 447.420 ;
        RECT 2.400 445.420 2497.200 446.780 ;
        RECT 2.400 425.660 2497.600 445.420 ;
        RECT 2.800 424.300 2497.600 425.660 ;
        RECT 2.800 423.660 2497.200 424.300 ;
        RECT 2.400 422.300 2497.200 423.660 ;
        RECT 2.400 403.900 2497.600 422.300 ;
        RECT 2.800 402.540 2497.600 403.900 ;
        RECT 2.800 401.900 2497.200 402.540 ;
        RECT 2.400 400.540 2497.200 401.900 ;
        RECT 2.400 380.780 2497.600 400.540 ;
        RECT 2.800 379.420 2497.600 380.780 ;
        RECT 2.800 378.780 2497.200 379.420 ;
        RECT 2.400 377.420 2497.200 378.780 ;
        RECT 2.400 359.020 2497.600 377.420 ;
        RECT 2.800 357.660 2497.600 359.020 ;
        RECT 2.800 357.020 2497.200 357.660 ;
        RECT 2.400 355.660 2497.200 357.020 ;
        RECT 2.400 335.900 2497.600 355.660 ;
        RECT 2.800 333.900 2497.200 335.900 ;
        RECT 2.400 314.140 2497.600 333.900 ;
        RECT 2.800 312.780 2497.600 314.140 ;
        RECT 2.800 312.140 2497.200 312.780 ;
        RECT 2.400 310.780 2497.200 312.140 ;
        RECT 2.400 291.020 2497.600 310.780 ;
        RECT 2.800 289.020 2497.200 291.020 ;
        RECT 2.400 269.260 2497.600 289.020 ;
        RECT 2.800 267.900 2497.600 269.260 ;
        RECT 2.800 267.260 2497.200 267.900 ;
        RECT 2.400 265.900 2497.200 267.260 ;
        RECT 2.400 247.500 2497.600 265.900 ;
        RECT 2.800 246.140 2497.600 247.500 ;
        RECT 2.800 245.500 2497.200 246.140 ;
        RECT 2.400 244.140 2497.200 245.500 ;
        RECT 2.400 224.380 2497.600 244.140 ;
        RECT 2.800 223.020 2497.600 224.380 ;
        RECT 2.800 222.380 2497.200 223.020 ;
        RECT 2.400 221.020 2497.200 222.380 ;
        RECT 2.400 202.620 2497.600 221.020 ;
        RECT 2.800 201.260 2497.600 202.620 ;
        RECT 2.800 200.620 2497.200 201.260 ;
        RECT 2.400 199.260 2497.200 200.620 ;
        RECT 2.400 179.500 2497.600 199.260 ;
        RECT 2.800 178.140 2497.600 179.500 ;
        RECT 2.800 177.500 2497.200 178.140 ;
        RECT 2.400 176.140 2497.200 177.500 ;
        RECT 2.400 157.740 2497.600 176.140 ;
        RECT 2.800 156.380 2497.600 157.740 ;
        RECT 2.800 155.740 2497.200 156.380 ;
        RECT 2.400 154.380 2497.200 155.740 ;
        RECT 2.400 134.620 2497.600 154.380 ;
        RECT 2.800 133.260 2497.600 134.620 ;
        RECT 2.800 132.620 2497.200 133.260 ;
        RECT 2.400 131.260 2497.200 132.620 ;
        RECT 2.400 112.860 2497.600 131.260 ;
        RECT 2.800 111.500 2497.600 112.860 ;
        RECT 2.800 110.860 2497.200 111.500 ;
        RECT 2.400 109.500 2497.200 110.860 ;
        RECT 2.400 89.740 2497.600 109.500 ;
        RECT 2.800 88.380 2497.600 89.740 ;
        RECT 2.800 87.740 2497.200 88.380 ;
        RECT 2.400 86.380 2497.200 87.740 ;
        RECT 2.400 67.980 2497.600 86.380 ;
        RECT 2.800 66.620 2497.600 67.980 ;
        RECT 2.800 65.980 2497.200 66.620 ;
        RECT 2.400 64.620 2497.200 65.980 ;
        RECT 2.400 44.860 2497.600 64.620 ;
        RECT 2.800 42.860 2497.200 44.860 ;
        RECT 2.400 23.100 2497.600 42.860 ;
        RECT 2.800 21.740 2497.600 23.100 ;
        RECT 2.800 21.100 2497.200 21.740 ;
        RECT 2.400 19.740 2497.200 21.100 ;
        RECT 2.400 15.135 2497.600 19.740 ;
      LAYER met4 ;
        RECT 71.040 15.135 1531.840 3084.305 ;
  END
END top
END LIBRARY

