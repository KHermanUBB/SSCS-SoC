VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.710 -4.800 2602.270 2.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1362.460 2924.800 1363.660 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 851.100 2.400 852.300 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.710 3517.600 1130.270 3524.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2189.340 2924.800 2190.540 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 3517.600 990.430 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 411.820 2.400 413.020 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3350.780 2924.800 3351.980 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1316.220 2.400 1317.420 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.190 3517.600 1216.750 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.750 -4.800 244.310 2.400 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.470 3517.600 903.030 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.310 3517.600 1042.870 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 360.140 2.400 361.340 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 980.300 2.400 981.500 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2525.260 2924.800 2526.460 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.630 3517.600 326.190 3524.800 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.390 3517.600 1915.950 3524.800 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.910 3517.600 955.470 3524.800 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 153.420 2.400 154.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.430 3517.600 1443.990 3524.800 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3201.180 2.400 3202.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.230 -4.800 1135.790 2.400 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1135.340 2.400 1136.540 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.230 3517.600 2055.790 3524.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.030 3517.600 1793.590 3524.800 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.110 -4.800 803.670 2.400 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2215.180 2924.800 2216.380 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1342.060 2.400 1343.260 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.870 -4.800 2462.430 2.400 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1367.900 2.400 1369.100 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.990 3517.600 2771.550 3524.800 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 123.500 2924.800 124.700 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1930.940 2924.800 1932.140 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2167.580 2.400 2168.780 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.350 3517.600 1513.910 3524.800 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2529.340 2.400 2530.540 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1026.540 2924.800 1027.740 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 949.020 2924.800 950.220 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.990 3517.600 1828.550 3524.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.750 3517.600 1164.310 3524.800 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.350 -4.800 1973.910 2.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.710 3517.600 693.270 3524.800 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1052.380 2924.800 1053.580 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.030 -4.800 1816.590 2.400 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 3517.600 238.790 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 3517.600 291.230 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1187.020 2.400 1188.220 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.190 3517.600 710.750 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.710 3517.600 2073.270 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 696.060 2.400 697.260 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1233.260 2924.800 1234.460 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3479.980 2924.800 3481.180 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3046.140 2.400 3047.340 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.390 3517.600 535.950 3524.800 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 50.060 2.400 51.260 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.950 3517.600 1863.510 3524.800 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2499.420 2924.800 2500.620 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2989.020 2924.800 2990.220 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.710 -4.800 1659.270 2.400 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3433.740 2.400 3434.940 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.350 3517.600 570.910 3524.800 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.110 3517.600 343.670 3524.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.670 3517.600 728.230 3524.800 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2115.900 2.400 2117.100 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.750 -4.800 1187.310 2.400 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2865.260 2.400 2866.460 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.470 3517.600 2283.030 3524.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1057.820 2.400 1059.020 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 3517.600 2160.670 3524.800 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2823.430 3517.600 2823.990 3524.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2761.900 2.400 2763.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.430 3517.600 500.990 3524.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 3517.600 203.830 3524.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.510 3517.600 2754.070 3524.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1779.980 2.400 1781.180 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3247.420 2924.800 3248.620 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1264.540 2.400 1265.740 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.630 -4.800 349.190 2.400 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2653.100 2924.800 2654.300 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 536.940 2924.800 538.140 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2163.500 2924.800 2164.700 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3118.220 2924.800 3119.420 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2678.940 2924.800 2680.140 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.670 -4.800 314.230 2.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.270 -4.800 2043.830 2.400 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 3517.600 168.870 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2531.790 -4.800 2532.350 2.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.910 -4.800 1484.470 2.400 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 71.820 2924.800 73.020 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2658.540 2.400 2659.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.630 3517.600 763.190 3524.800 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.630 -4.800 2672.190 2.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1801.740 2924.800 1802.940 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.310 -4.800 628.870 2.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2805.950 3517.600 2806.510 3524.800 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.070 -4.800 838.630 2.400 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3066.540 2924.800 3067.740 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2409.430 -4.800 2409.990 2.400 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2576.940 2924.800 2578.140 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2893.350 3517.600 2893.910 3524.800 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2266.860 2924.800 2268.060 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.150 3517.600 745.710 3524.800 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2391.950 -4.800 2392.510 2.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1909.180 2.400 1910.380 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 20.140 2924.800 21.340 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2060.140 2924.800 2061.340 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.270 3517.600 1583.830 3524.800 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 902.780 2.400 903.980 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.070 3517.600 1321.630 3524.800 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 3517.600 186.350 3524.800 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.550 -4.800 856.110 2.400 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1207.420 2924.800 1208.620 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 3517.600 2352.030 3524.800 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1620.860 2924.800 1622.060 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 743.660 2924.800 744.860 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.470 3517.600 1409.030 3524.800 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.750 3517.600 658.310 3524.800 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3195.740 2924.800 3196.940 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2942.780 2.400 2943.980 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2085.980 2924.800 2087.180 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 45.980 2924.800 47.180 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.150 3517.600 1688.710 3524.800 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 666.140 2924.800 667.340 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.630 3517.600 2143.190 3524.800 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3020.300 2.400 3021.500 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 -4.800 86.990 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2111.820 2924.800 2113.020 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3071.980 2.400 3073.180 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 252.700 2924.800 253.900 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.550 3517.600 2213.110 3524.800 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.790 -4.800 646.350 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.190 -4.800 1170.750 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.590 3517.600 1304.150 3524.800 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.430 3517.600 2386.990 3524.800 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1982.620 2924.800 1983.820 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2813.580 2.400 2814.780 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.750 3517.600 2038.310 3524.800 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2584.230 -4.800 2584.790 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 3517.600 361.150 3524.800 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2706.590 -4.800 2707.150 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.470 3517.600 466.030 3524.800 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1006.140 2.400 1007.340 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.790 -4.800 2026.350 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2090.060 2.400 2091.260 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1754.140 2.400 1755.340 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.990 -4.800 2357.550 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2447.740 2924.800 2448.940 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 618.540 2.400 619.740 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1284.940 2924.800 1286.140 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1600.460 2.400 1601.660 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2911.500 2924.800 2912.700 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.990 3517.600 2265.550 3524.800 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.270 -4.800 663.830 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.190 3517.600 273.750 3524.800 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 127.580 2.400 128.780 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.590 -4.800 1764.150 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1698.380 2924.800 1699.580 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 407.740 2924.800 408.940 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2581.020 2.400 2582.220 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2756.460 2924.800 2757.660 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 282.620 2.400 283.820 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1956.780 2924.800 1957.980 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.430 -4.800 1903.990 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.190 -4.800 2113.750 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.710 3517.600 1199.270 3524.800 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.390 -4.800 1938.950 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.270 -4.800 1100.830 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.910 3517.600 1461.470 3524.800 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3252.860 2.400 3254.060 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 3517.600 2334.550 3524.800 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2840.910 3517.600 2841.470 3524.800 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1336.620 2924.800 1337.820 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 -4.800 52.030 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2012.540 2.400 2013.740 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.910 -4.800 541.470 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1414.140 2924.800 1415.340 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2628.620 2924.800 2629.820 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.230 3517.600 1112.790 3524.800 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 670.220 2.400 671.420 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2141.740 2.400 2142.940 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.070 -4.800 1781.630 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.150 3517.600 2125.710 3524.800 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.430 -4.800 523.990 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.470 -4.800 926.030 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 75.900 2.400 77.100 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 3517.600 256.270 3524.800 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2788.470 3517.600 2789.030 3524.800 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 381.900 2924.800 383.100 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.150 -4.800 331.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.670 -4.800 1257.230 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 -4.800 17.070 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.830 -4.800 1991.390 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.350 3517.600 2456.910 3524.800 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.950 -4.800 2323.510 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1652.140 2.400 1653.340 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 3517.600 431.070 3524.800 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.390 -4.800 558.950 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 588.620 2924.800 589.820 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2193.420 2.400 2194.620 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3299.100 2924.800 3300.300 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2305.470 -4.800 2306.030 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 3517.600 98.950 3524.800 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 3517.600 1339.110 3524.800 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 954.460 2.400 955.660 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2473.580 2924.800 2474.780 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1181.580 2924.800 1182.780 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 614.460 2924.800 615.660 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 356.060 2924.800 357.260 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.990 3517.600 885.550 3524.800 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2636.670 -4.800 2637.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.110 -4.800 1309.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.830 -4.800 1048.390 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.630 -4.800 1292.190 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2137.660 2924.800 2138.860 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2730.620 2924.800 2731.820 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 717.820 2924.800 719.020 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 847.020 2924.800 848.220 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.110 -4.800 2183.670 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 872.860 2924.800 874.060 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1729.660 2.400 1730.860 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 24.220 2.400 25.420 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.110 3517.600 1286.670 3524.800 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2396.060 2924.800 2397.260 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1960.860 2.400 1962.060 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2374.300 2.400 2375.500 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.190 3517.600 1147.750 3524.800 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.030 3517.600 850.590 3524.800 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1775.550 3517.600 1776.110 3524.800 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.150 3517.600 308.710 3524.800 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2724.070 -4.800 2724.630 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.950 -4.800 943.510 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.310 -4.800 1065.870 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1393.740 2.400 1394.940 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3407.900 2.400 3409.100 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1465.820 2924.800 1467.020 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2632.700 2.400 2633.900 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.990 -4.800 471.550 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2451.820 2.400 2453.020 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2718.550 3517.600 2719.110 3524.800 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3382.060 2.400 3383.260 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 334.300 2.400 335.500 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1078.220 2924.800 1079.420 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1750.060 2924.800 1751.260 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1238.700 2.400 1239.900 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.550 3517.600 833.110 3524.800 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3097.820 2.400 3099.020 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.230 3517.600 1618.790 3524.800 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.470 3517.600 1846.030 3524.800 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.550 -4.800 419.110 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.070 3517.600 2195.630 3524.800 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2666.110 3517.600 2666.670 3524.800 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 308.460 2.400 309.660 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 3517.600 1356.590 3524.800 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3040.700 2924.800 3041.900 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 511.100 2924.800 512.300 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 928.620 2.400 929.820 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.870 -4.800 1013.430 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1419.580 2.400 1420.780 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.030 -4.800 2759.590 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.230 3517.600 675.790 3524.800 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.070 3517.600 2701.630 3524.800 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1290.380 2.400 1291.580 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2426.910 -4.800 2427.470 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.350 -4.800 1536.910 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2348.460 2.400 2349.660 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3092.380 2924.800 3093.580 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1388.300 2924.800 1389.500 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1522.940 2.400 1524.140 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1569.180 2924.800 1570.380 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.990 3517.600 448.550 3524.800 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 304.380 2924.800 305.580 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2503.500 2.400 2504.700 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 3517.600 413.590 3524.800 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3402.460 2924.800 3403.660 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 799.420 2.400 800.620 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.310 3517.600 1985.870 3524.800 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1104.060 2924.800 1105.260 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.110 3517.600 1723.670 3524.800 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 773.580 2.400 774.780 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1439.980 2924.800 1441.180 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.430 3517.600 63.990 3524.800 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 201.020 2924.800 202.220 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.190 -4.800 1239.750 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1161.180 2.400 1162.380 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.590 3517.600 798.150 3524.800 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 3517.600 1758.630 3524.800 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.750 -4.800 2567.310 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.190 3517.600 2596.750 3524.800 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2916.940 2.400 2918.140 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1857.500 2.400 1858.700 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.950 3517.600 2369.510 3524.800 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 691.980 2924.800 693.180 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.150 3517.600 1251.710 3524.800 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2477.660 2.400 2478.860 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.790 3517.600 1060.350 3524.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.390 3517.600 972.950 3524.800 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.550 -4.800 2236.110 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2741.550 -4.800 2742.110 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.870 3517.600 2876.430 3524.800 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.230 3517.600 1181.790 3524.800 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 463.500 2.400 464.700 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.310 -4.800 191.870 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1831.660 2.400 1832.860 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2219.260 2.400 2220.460 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.590 -4.800 821.150 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2968.620 2.400 2969.820 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1595.020 2924.800 1596.220 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2400.140 2.400 2401.340 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1491.660 2924.800 1492.860 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 205.100 2.400 206.300 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.510 -4.800 1397.070 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.030 3517.600 2736.590 3524.800 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.950 3517.600 2300.510 3524.800 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 3517.600 1531.390 3524.800 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.110 -4.800 366.670 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3330.380 2.400 3331.580 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1724.220 2924.800 1725.420 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 485.260 2924.800 486.460 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 149.340 2924.800 150.540 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.150 -4.800 1274.710 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.950 -4.800 1886.510 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2648.630 3517.600 2649.190 3524.800 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.950 -4.800 1449.510 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.630 3517.600 1269.190 3524.800 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 3517.600 116.430 3524.800 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.710 -4.800 716.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.790 3517.600 1566.350 3524.800 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.350 -4.800 2916.910 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.310 -4.800 2514.870 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 459.420 2924.800 460.620 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 278.540 2924.800 279.740 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 3517.600 46.510 3524.800 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 489.340 2.400 490.540 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.070 3517.600 815.630 3524.800 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.630 -4.800 2166.190 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.790 3517.600 623.350 3524.800 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 721.900 2.400 723.100 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.150 -4.800 2654.710 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1646.700 2924.800 1647.900 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.630 3517.600 1706.190 3524.800 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.670 -4.800 1694.230 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.710 3517.600 1636.270 3524.800 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.190 3517.600 1653.750 3524.800 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.310 -4.800 2008.870 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.030 -4.800 2253.590 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 3517.600 2509.350 3524.800 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.510 3517.600 1374.070 3524.800 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.950 3517.600 483.510 3524.800 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.870 3517.600 2439.430 3524.800 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2689.110 -4.800 2689.670 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.230 -4.800 1204.790 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.990 -4.800 1414.550 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3454.140 2924.800 3455.340 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3278.700 2.400 3279.900 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.310 3517.600 2491.870 3524.800 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.750 -4.800 681.310 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1879.260 2924.800 1880.460 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.390 3517.600 1478.950 3524.800 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2858.390 3517.600 2858.950 3524.800 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1827.580 2924.800 1828.780 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.790 3517.600 2003.350 3524.800 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.430 3517.600 2317.990 3524.800 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.790 -4.800 1083.350 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2602.780 2924.800 2603.980 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.870 -4.800 1956.430 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2038.380 2.400 2039.580 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.950 -4.800 506.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 3517.600 1811.070 3524.800 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.830 -4.800 1554.390 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.030 -4.800 1379.590 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3324.940 2924.800 3326.140 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1155.740 2924.800 1156.940 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1883.340 2.400 1884.540 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1853.420 2924.800 1854.620 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.150 -4.800 1711.710 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.430 -4.800 960.990 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2839.420 2.400 2840.620 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2859.820 2924.800 2861.020 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2270.940 2.400 2272.140 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2684.380 2.400 2685.580 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.590 -4.800 2201.150 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 640.300 2924.800 641.500 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2318.540 2924.800 2319.740 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 644.380 2.400 645.580 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 541.020 2.400 542.220 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.470 -4.800 1432.030 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.150 -4.800 768.710 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 330.220 2924.800 331.420 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.630 -4.800 786.190 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 226.860 2924.800 228.060 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3273.260 2924.800 3274.460 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1259.100 2924.800 1260.300 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 -4.800 279.270 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1212.860 2.400 1214.060 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.470 -4.800 1869.030 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2578.710 3517.600 2579.270 3524.800 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1775.900 2924.800 1777.100 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 3517.600 2911.390 3524.800 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.670 3517.600 2614.230 3524.800 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 179.260 2.400 180.460 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1805.820 2.400 1807.020 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 3517.600 1007.910 3524.800 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.510 -4.800 891.070 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.870 3517.600 553.430 3524.800 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 898.700 2924.800 899.900 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.100 2924.800 1906.300 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 515.180 2.400 516.380 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.750 -4.800 2061.310 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2808.140 2924.800 2809.340 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2606.860 2.400 2608.060 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2683.590 3517.600 2684.150 3524.800 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3356.220 2.400 3357.420 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.070 3517.600 378.630 3524.800 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3304.540 2.400 3305.740 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2846.430 -4.800 2846.990 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.470 -4.800 489.030 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.190 -4.800 733.750 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.270 -4.800 2549.830 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 821.180 2924.800 822.380 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2833.980 2924.800 2835.180 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2710.220 2.400 2711.420 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.870 3517.600 1496.430 3524.800 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.270 3517.600 1077.830 3524.800 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1935.020 2.400 1936.220 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3221.580 2924.800 3222.780 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2891.100 2.400 2892.300 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.950 3517.600 920.510 3524.800 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 566.860 2.400 568.060 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2782.300 2924.800 2783.500 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 3517.600 2108.230 3524.800 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 3517.600 81.470 3524.800 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2403.910 3517.600 2404.470 3524.800 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.750 3517.600 2544.310 3524.800 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2561.230 3517.600 2561.790 3524.800 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.790 -4.800 1589.350 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.670 3517.600 1671.230 3524.800 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 -4.800 104.470 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 -4.800 34.550 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2374.470 -4.800 2375.030 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1626.300 2.400 1627.500 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 433.580 2924.800 434.780 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2064.220 2.400 2065.420 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2736.060 2.400 2737.260 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 3517.600 151.390 3524.800 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1703.820 2.400 1705.020 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1445.420 2.400 1446.620 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1109.500 2.400 1110.700 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.750 3517.600 1601.310 3524.800 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.390 -4.800 2444.950 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.710 -4.800 1153.270 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3175.340 2.400 3176.540 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2344.380 2924.800 2345.580 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3169.900 2924.800 3171.100 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2296.780 2.400 2297.980 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2787.740 2.400 2788.940 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 97.660 2924.800 98.860 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2963.180 2924.800 2964.380 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.670 3517.600 1234.230 3524.800 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2421.900 2924.800 2423.100 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.990 -4.800 2288.550 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 562.780 2924.800 563.980 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.830 3517.600 1025.390 3524.800 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.510 -4.800 2777.070 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 3517.600 11.550 3524.800 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.590 -4.800 384.150 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1497.100 2.400 1498.300 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.190 -4.800 1676.750 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2937.340 2924.800 2938.540 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.670 -4.800 751.230 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2811.470 -4.800 2812.030 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.750 3517.600 221.310 3524.800 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.910 3517.600 1898.470 3524.800 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 592.700 2.400 593.900 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 3517.600 133.910 3524.800 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.550 3517.600 396.110 3524.800 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 795.340 2924.800 796.540 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3484.060 2.400 3485.260 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1083.660 2.400 1084.860 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.990 3517.600 1391.550 3524.800 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.110 3517.600 780.670 3524.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2994.460 2.400 2995.660 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 -4.800 261.790 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2322.620 2.400 2323.820 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3144.060 2924.800 3145.260 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2885.660 2924.800 2886.860 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.990 -4.800 1851.550 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 256.780 2.400 257.980 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1310.780 2924.800 1311.980 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2793.990 -4.800 2794.550 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.950 3517.600 1426.510 3524.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.510 3517.600 2248.070 3524.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.230 -4.800 1641.790 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.430 -4.800 2340.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 923.180 2924.800 924.380 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3459.580 2.400 3460.780 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.310 -4.800 1571.870 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 -4.800 296.750 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 3517.600 605.870 3524.800 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2370.220 2924.800 2371.420 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.150 3517.600 2631.710 3524.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.750 -4.800 1118.310 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.870 3517.600 1933.430 3524.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1672.540 2924.800 1673.740 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.070 -4.800 2218.630 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.430 3517.600 1880.990 3524.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.990 -4.800 908.550 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 -4.800 139.430 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.950 -4.800 2829.510 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1000.700 2924.800 1001.900 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.270 3517.600 640.830 3524.800 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3505.820 2924.800 3507.020 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2245.100 2.400 2246.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2555.180 2.400 2556.380 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 385.980 2.400 387.180 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.830 -4.800 611.390 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2008.460 2924.800 2009.660 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.270 -4.800 1606.830 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.590 3517.600 1741.150 3524.800 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2421.390 3517.600 2421.950 3524.800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3509.900 2.400 3511.100 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.030 -4.800 436.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2292.700 2924.800 2293.900 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.270 3517.600 2526.830 3524.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1677.980 2.400 1679.180 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3014.860 2924.800 3016.060 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1129.900 2924.800 1131.100 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 101.740 2.400 102.940 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.030 3517.600 2230.590 3524.800 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 3517.600 588.390 3524.800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.030 -4.800 873.590 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2241.020 2924.800 2242.220 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.510 -4.800 2271.070 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 974.860 2924.800 976.060 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1548.780 2.400 1549.980 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.910 -4.800 2864.470 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.510 -4.800 454.070 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.550 -4.800 1362.110 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1517.500 2924.800 1518.700 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 3517.600 2178.150 3524.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3376.620 2924.800 3377.820 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.270 -4.800 226.830 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2034.300 2924.800 2035.500 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 -4.800 69.510 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3428.300 2924.800 3429.500 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.190 3517.600 2090.750 3524.800 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 175.180 2924.800 176.380 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 437.660 2.400 438.860 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 747.740 2.400 748.940 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 876.940 2.400 878.140 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.510 -4.800 1834.070 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 -4.800 0.510 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1574.620 2.400 1575.820 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3149.500 2.400 3150.700 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.510 3517.600 868.070 3524.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1031.980 2.400 1033.180 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 -4.800 209.350 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.310 3517.600 1548.870 3524.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.430 3517.600 937.990 3524.800 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.430 -4.800 1466.990 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2020.270 3517.600 2020.830 3524.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 769.500 2924.800 770.700 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2425.980 2.400 2427.180 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2704.780 2924.800 2705.980 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.350 -4.800 593.910 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.350 -4.800 1030.910 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 230.940 2.400 232.140 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.750 -4.800 1624.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.830 3517.600 1968.390 3524.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.350 3517.600 1950.910 3524.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 3517.600 29.030 3524.800 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.910 3517.600 518.470 3524.800 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.910 -4.800 1921.470 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 825.260 2.400 826.460 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3227.020 2.400 3228.220 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1543.340 2924.800 1544.540 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 7.820 17.085 2912.115 3503.445 ;
      LAYER met1 ;
        RECT 0.070 13.980 2916.790 3515.220 ;
      LAYER met2 ;
        RECT 0.100 3517.320 10.710 3518.050 ;
        RECT 11.830 3517.320 28.190 3518.050 ;
        RECT 29.310 3517.320 45.670 3518.050 ;
        RECT 46.790 3517.320 63.150 3518.050 ;
        RECT 64.270 3517.320 80.630 3518.050 ;
        RECT 81.750 3517.320 98.110 3518.050 ;
        RECT 99.230 3517.320 115.590 3518.050 ;
        RECT 116.710 3517.320 133.070 3518.050 ;
        RECT 134.190 3517.320 150.550 3518.050 ;
        RECT 151.670 3517.320 168.030 3518.050 ;
        RECT 169.150 3517.320 185.510 3518.050 ;
        RECT 186.630 3517.320 202.990 3518.050 ;
        RECT 204.110 3517.320 220.470 3518.050 ;
        RECT 221.590 3517.320 237.950 3518.050 ;
        RECT 239.070 3517.320 255.430 3518.050 ;
        RECT 256.550 3517.320 272.910 3518.050 ;
        RECT 274.030 3517.320 290.390 3518.050 ;
        RECT 291.510 3517.320 307.870 3518.050 ;
        RECT 308.990 3517.320 325.350 3518.050 ;
        RECT 326.470 3517.320 342.830 3518.050 ;
        RECT 343.950 3517.320 360.310 3518.050 ;
        RECT 361.430 3517.320 377.790 3518.050 ;
        RECT 378.910 3517.320 395.270 3518.050 ;
        RECT 396.390 3517.320 412.750 3518.050 ;
        RECT 413.870 3517.320 430.230 3518.050 ;
        RECT 431.350 3517.320 447.710 3518.050 ;
        RECT 448.830 3517.320 465.190 3518.050 ;
        RECT 466.310 3517.320 482.670 3518.050 ;
        RECT 483.790 3517.320 500.150 3518.050 ;
        RECT 501.270 3517.320 517.630 3518.050 ;
        RECT 518.750 3517.320 535.110 3518.050 ;
        RECT 536.230 3517.320 552.590 3518.050 ;
        RECT 553.710 3517.320 570.070 3518.050 ;
        RECT 571.190 3517.320 587.550 3518.050 ;
        RECT 588.670 3517.320 605.030 3518.050 ;
        RECT 606.150 3517.320 622.510 3518.050 ;
        RECT 623.630 3517.320 639.990 3518.050 ;
        RECT 641.110 3517.320 657.470 3518.050 ;
        RECT 658.590 3517.320 674.950 3518.050 ;
        RECT 676.070 3517.320 692.430 3518.050 ;
        RECT 693.550 3517.320 709.910 3518.050 ;
        RECT 711.030 3517.320 727.390 3518.050 ;
        RECT 728.510 3517.320 744.870 3518.050 ;
        RECT 745.990 3517.320 762.350 3518.050 ;
        RECT 763.470 3517.320 779.830 3518.050 ;
        RECT 780.950 3517.320 797.310 3518.050 ;
        RECT 798.430 3517.320 814.790 3518.050 ;
        RECT 815.910 3517.320 832.270 3518.050 ;
        RECT 833.390 3517.320 849.750 3518.050 ;
        RECT 850.870 3517.320 867.230 3518.050 ;
        RECT 868.350 3517.320 884.710 3518.050 ;
        RECT 885.830 3517.320 902.190 3518.050 ;
        RECT 903.310 3517.320 919.670 3518.050 ;
        RECT 920.790 3517.320 937.150 3518.050 ;
        RECT 938.270 3517.320 954.630 3518.050 ;
        RECT 955.750 3517.320 972.110 3518.050 ;
        RECT 973.230 3517.320 989.590 3518.050 ;
        RECT 990.710 3517.320 1007.070 3518.050 ;
        RECT 1008.190 3517.320 1024.550 3518.050 ;
        RECT 1025.670 3517.320 1042.030 3518.050 ;
        RECT 1043.150 3517.320 1059.510 3518.050 ;
        RECT 1060.630 3517.320 1076.990 3518.050 ;
        RECT 1078.110 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1111.950 3518.050 ;
        RECT 1113.070 3517.320 1129.430 3518.050 ;
        RECT 1130.550 3517.320 1146.910 3518.050 ;
        RECT 1148.030 3517.320 1163.470 3518.050 ;
        RECT 1164.590 3517.320 1180.950 3518.050 ;
        RECT 1182.070 3517.320 1198.430 3518.050 ;
        RECT 1199.550 3517.320 1215.910 3518.050 ;
        RECT 1217.030 3517.320 1233.390 3518.050 ;
        RECT 1234.510 3517.320 1250.870 3518.050 ;
        RECT 1251.990 3517.320 1268.350 3518.050 ;
        RECT 1269.470 3517.320 1285.830 3518.050 ;
        RECT 1286.950 3517.320 1303.310 3518.050 ;
        RECT 1304.430 3517.320 1320.790 3518.050 ;
        RECT 1321.910 3517.320 1338.270 3518.050 ;
        RECT 1339.390 3517.320 1355.750 3518.050 ;
        RECT 1356.870 3517.320 1373.230 3518.050 ;
        RECT 1374.350 3517.320 1390.710 3518.050 ;
        RECT 1391.830 3517.320 1408.190 3518.050 ;
        RECT 1409.310 3517.320 1425.670 3518.050 ;
        RECT 1426.790 3517.320 1443.150 3518.050 ;
        RECT 1444.270 3517.320 1460.630 3518.050 ;
        RECT 1461.750 3517.320 1478.110 3518.050 ;
        RECT 1479.230 3517.320 1495.590 3518.050 ;
        RECT 1496.710 3517.320 1513.070 3518.050 ;
        RECT 1514.190 3517.320 1530.550 3518.050 ;
        RECT 1531.670 3517.320 1548.030 3518.050 ;
        RECT 1549.150 3517.320 1565.510 3518.050 ;
        RECT 1566.630 3517.320 1582.990 3518.050 ;
        RECT 1584.110 3517.320 1600.470 3518.050 ;
        RECT 1601.590 3517.320 1617.950 3518.050 ;
        RECT 1619.070 3517.320 1635.430 3518.050 ;
        RECT 1636.550 3517.320 1652.910 3518.050 ;
        RECT 1654.030 3517.320 1670.390 3518.050 ;
        RECT 1671.510 3517.320 1687.870 3518.050 ;
        RECT 1688.990 3517.320 1705.350 3518.050 ;
        RECT 1706.470 3517.320 1722.830 3518.050 ;
        RECT 1723.950 3517.320 1740.310 3518.050 ;
        RECT 1741.430 3517.320 1757.790 3518.050 ;
        RECT 1758.910 3517.320 1775.270 3518.050 ;
        RECT 1776.390 3517.320 1792.750 3518.050 ;
        RECT 1793.870 3517.320 1810.230 3518.050 ;
        RECT 1811.350 3517.320 1827.710 3518.050 ;
        RECT 1828.830 3517.320 1845.190 3518.050 ;
        RECT 1846.310 3517.320 1862.670 3518.050 ;
        RECT 1863.790 3517.320 1880.150 3518.050 ;
        RECT 1881.270 3517.320 1897.630 3518.050 ;
        RECT 1898.750 3517.320 1915.110 3518.050 ;
        RECT 1916.230 3517.320 1932.590 3518.050 ;
        RECT 1933.710 3517.320 1950.070 3518.050 ;
        RECT 1951.190 3517.320 1967.550 3518.050 ;
        RECT 1968.670 3517.320 1985.030 3518.050 ;
        RECT 1986.150 3517.320 2002.510 3518.050 ;
        RECT 2003.630 3517.320 2019.990 3518.050 ;
        RECT 2021.110 3517.320 2037.470 3518.050 ;
        RECT 2038.590 3517.320 2054.950 3518.050 ;
        RECT 2056.070 3517.320 2072.430 3518.050 ;
        RECT 2073.550 3517.320 2089.910 3518.050 ;
        RECT 2091.030 3517.320 2107.390 3518.050 ;
        RECT 2108.510 3517.320 2124.870 3518.050 ;
        RECT 2125.990 3517.320 2142.350 3518.050 ;
        RECT 2143.470 3517.320 2159.830 3518.050 ;
        RECT 2160.950 3517.320 2177.310 3518.050 ;
        RECT 2178.430 3517.320 2194.790 3518.050 ;
        RECT 2195.910 3517.320 2212.270 3518.050 ;
        RECT 2213.390 3517.320 2229.750 3518.050 ;
        RECT 2230.870 3517.320 2247.230 3518.050 ;
        RECT 2248.350 3517.320 2264.710 3518.050 ;
        RECT 2265.830 3517.320 2282.190 3518.050 ;
        RECT 2283.310 3517.320 2299.670 3518.050 ;
        RECT 2300.790 3517.320 2317.150 3518.050 ;
        RECT 2318.270 3517.320 2333.710 3518.050 ;
        RECT 2334.830 3517.320 2351.190 3518.050 ;
        RECT 2352.310 3517.320 2368.670 3518.050 ;
        RECT 2369.790 3517.320 2386.150 3518.050 ;
        RECT 2387.270 3517.320 2403.630 3518.050 ;
        RECT 2404.750 3517.320 2421.110 3518.050 ;
        RECT 2422.230 3517.320 2438.590 3518.050 ;
        RECT 2439.710 3517.320 2456.070 3518.050 ;
        RECT 2457.190 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2491.030 3518.050 ;
        RECT 2492.150 3517.320 2508.510 3518.050 ;
        RECT 2509.630 3517.320 2525.990 3518.050 ;
        RECT 2527.110 3517.320 2543.470 3518.050 ;
        RECT 2544.590 3517.320 2560.950 3518.050 ;
        RECT 2562.070 3517.320 2578.430 3518.050 ;
        RECT 2579.550 3517.320 2595.910 3518.050 ;
        RECT 2597.030 3517.320 2613.390 3518.050 ;
        RECT 2614.510 3517.320 2630.870 3518.050 ;
        RECT 2631.990 3517.320 2648.350 3518.050 ;
        RECT 2649.470 3517.320 2665.830 3518.050 ;
        RECT 2666.950 3517.320 2683.310 3518.050 ;
        RECT 2684.430 3517.320 2700.790 3518.050 ;
        RECT 2701.910 3517.320 2718.270 3518.050 ;
        RECT 2719.390 3517.320 2735.750 3518.050 ;
        RECT 2736.870 3517.320 2753.230 3518.050 ;
        RECT 2754.350 3517.320 2770.710 3518.050 ;
        RECT 2771.830 3517.320 2788.190 3518.050 ;
        RECT 2789.310 3517.320 2805.670 3518.050 ;
        RECT 2806.790 3517.320 2823.150 3518.050 ;
        RECT 2824.270 3517.320 2840.630 3518.050 ;
        RECT 2841.750 3517.320 2858.110 3518.050 ;
        RECT 2859.230 3517.320 2875.590 3518.050 ;
        RECT 2876.710 3517.320 2893.070 3518.050 ;
        RECT 2894.190 3517.320 2910.550 3518.050 ;
        RECT 2911.670 3517.320 2916.760 3518.050 ;
        RECT 0.100 2.680 2916.760 3517.320 ;
        RECT 0.790 2.310 16.230 2.680 ;
        RECT 17.350 2.310 33.710 2.680 ;
        RECT 34.830 2.310 51.190 2.680 ;
        RECT 52.310 2.310 68.670 2.680 ;
        RECT 69.790 2.310 86.150 2.680 ;
        RECT 87.270 2.310 103.630 2.680 ;
        RECT 104.750 2.310 121.110 2.680 ;
        RECT 122.230 2.310 138.590 2.680 ;
        RECT 139.710 2.310 156.070 2.680 ;
        RECT 157.190 2.310 173.550 2.680 ;
        RECT 174.670 2.310 191.030 2.680 ;
        RECT 192.150 2.310 208.510 2.680 ;
        RECT 209.630 2.310 225.990 2.680 ;
        RECT 227.110 2.310 243.470 2.680 ;
        RECT 244.590 2.310 260.950 2.680 ;
        RECT 262.070 2.310 278.430 2.680 ;
        RECT 279.550 2.310 295.910 2.680 ;
        RECT 297.030 2.310 313.390 2.680 ;
        RECT 314.510 2.310 330.870 2.680 ;
        RECT 331.990 2.310 348.350 2.680 ;
        RECT 349.470 2.310 365.830 2.680 ;
        RECT 366.950 2.310 383.310 2.680 ;
        RECT 384.430 2.310 400.790 2.680 ;
        RECT 401.910 2.310 418.270 2.680 ;
        RECT 419.390 2.310 435.750 2.680 ;
        RECT 436.870 2.310 453.230 2.680 ;
        RECT 454.350 2.310 470.710 2.680 ;
        RECT 471.830 2.310 488.190 2.680 ;
        RECT 489.310 2.310 505.670 2.680 ;
        RECT 506.790 2.310 523.150 2.680 ;
        RECT 524.270 2.310 540.630 2.680 ;
        RECT 541.750 2.310 558.110 2.680 ;
        RECT 559.230 2.310 575.590 2.680 ;
        RECT 576.710 2.310 593.070 2.680 ;
        RECT 594.190 2.310 610.550 2.680 ;
        RECT 611.670 2.310 628.030 2.680 ;
        RECT 629.150 2.310 645.510 2.680 ;
        RECT 646.630 2.310 662.990 2.680 ;
        RECT 664.110 2.310 680.470 2.680 ;
        RECT 681.590 2.310 697.950 2.680 ;
        RECT 699.070 2.310 715.430 2.680 ;
        RECT 716.550 2.310 732.910 2.680 ;
        RECT 734.030 2.310 750.390 2.680 ;
        RECT 751.510 2.310 767.870 2.680 ;
        RECT 768.990 2.310 785.350 2.680 ;
        RECT 786.470 2.310 802.830 2.680 ;
        RECT 803.950 2.310 820.310 2.680 ;
        RECT 821.430 2.310 837.790 2.680 ;
        RECT 838.910 2.310 855.270 2.680 ;
        RECT 856.390 2.310 872.750 2.680 ;
        RECT 873.870 2.310 890.230 2.680 ;
        RECT 891.350 2.310 907.710 2.680 ;
        RECT 908.830 2.310 925.190 2.680 ;
        RECT 926.310 2.310 942.670 2.680 ;
        RECT 943.790 2.310 960.150 2.680 ;
        RECT 961.270 2.310 977.630 2.680 ;
        RECT 978.750 2.310 995.110 2.680 ;
        RECT 996.230 2.310 1012.590 2.680 ;
        RECT 1013.710 2.310 1030.070 2.680 ;
        RECT 1031.190 2.310 1047.550 2.680 ;
        RECT 1048.670 2.310 1065.030 2.680 ;
        RECT 1066.150 2.310 1082.510 2.680 ;
        RECT 1083.630 2.310 1099.990 2.680 ;
        RECT 1101.110 2.310 1117.470 2.680 ;
        RECT 1118.590 2.310 1134.950 2.680 ;
        RECT 1136.070 2.310 1152.430 2.680 ;
        RECT 1153.550 2.310 1169.910 2.680 ;
        RECT 1171.030 2.310 1186.470 2.680 ;
        RECT 1187.590 2.310 1203.950 2.680 ;
        RECT 1205.070 2.310 1221.430 2.680 ;
        RECT 1222.550 2.310 1238.910 2.680 ;
        RECT 1240.030 2.310 1256.390 2.680 ;
        RECT 1257.510 2.310 1273.870 2.680 ;
        RECT 1274.990 2.310 1291.350 2.680 ;
        RECT 1292.470 2.310 1308.830 2.680 ;
        RECT 1309.950 2.310 1326.310 2.680 ;
        RECT 1327.430 2.310 1343.790 2.680 ;
        RECT 1344.910 2.310 1361.270 2.680 ;
        RECT 1362.390 2.310 1378.750 2.680 ;
        RECT 1379.870 2.310 1396.230 2.680 ;
        RECT 1397.350 2.310 1413.710 2.680 ;
        RECT 1414.830 2.310 1431.190 2.680 ;
        RECT 1432.310 2.310 1448.670 2.680 ;
        RECT 1449.790 2.310 1466.150 2.680 ;
        RECT 1467.270 2.310 1483.630 2.680 ;
        RECT 1484.750 2.310 1501.110 2.680 ;
        RECT 1502.230 2.310 1518.590 2.680 ;
        RECT 1519.710 2.310 1536.070 2.680 ;
        RECT 1537.190 2.310 1553.550 2.680 ;
        RECT 1554.670 2.310 1571.030 2.680 ;
        RECT 1572.150 2.310 1588.510 2.680 ;
        RECT 1589.630 2.310 1605.990 2.680 ;
        RECT 1607.110 2.310 1623.470 2.680 ;
        RECT 1624.590 2.310 1640.950 2.680 ;
        RECT 1642.070 2.310 1658.430 2.680 ;
        RECT 1659.550 2.310 1675.910 2.680 ;
        RECT 1677.030 2.310 1693.390 2.680 ;
        RECT 1694.510 2.310 1710.870 2.680 ;
        RECT 1711.990 2.310 1728.350 2.680 ;
        RECT 1729.470 2.310 1745.830 2.680 ;
        RECT 1746.950 2.310 1763.310 2.680 ;
        RECT 1764.430 2.310 1780.790 2.680 ;
        RECT 1781.910 2.310 1798.270 2.680 ;
        RECT 1799.390 2.310 1815.750 2.680 ;
        RECT 1816.870 2.310 1833.230 2.680 ;
        RECT 1834.350 2.310 1850.710 2.680 ;
        RECT 1851.830 2.310 1868.190 2.680 ;
        RECT 1869.310 2.310 1885.670 2.680 ;
        RECT 1886.790 2.310 1903.150 2.680 ;
        RECT 1904.270 2.310 1920.630 2.680 ;
        RECT 1921.750 2.310 1938.110 2.680 ;
        RECT 1939.230 2.310 1955.590 2.680 ;
        RECT 1956.710 2.310 1973.070 2.680 ;
        RECT 1974.190 2.310 1990.550 2.680 ;
        RECT 1991.670 2.310 2008.030 2.680 ;
        RECT 2009.150 2.310 2025.510 2.680 ;
        RECT 2026.630 2.310 2042.990 2.680 ;
        RECT 2044.110 2.310 2060.470 2.680 ;
        RECT 2061.590 2.310 2077.950 2.680 ;
        RECT 2079.070 2.310 2095.430 2.680 ;
        RECT 2096.550 2.310 2112.910 2.680 ;
        RECT 2114.030 2.310 2130.390 2.680 ;
        RECT 2131.510 2.310 2147.870 2.680 ;
        RECT 2148.990 2.310 2165.350 2.680 ;
        RECT 2166.470 2.310 2182.830 2.680 ;
        RECT 2183.950 2.310 2200.310 2.680 ;
        RECT 2201.430 2.310 2217.790 2.680 ;
        RECT 2218.910 2.310 2235.270 2.680 ;
        RECT 2236.390 2.310 2252.750 2.680 ;
        RECT 2253.870 2.310 2270.230 2.680 ;
        RECT 2271.350 2.310 2287.710 2.680 ;
        RECT 2288.830 2.310 2305.190 2.680 ;
        RECT 2306.310 2.310 2322.670 2.680 ;
        RECT 2323.790 2.310 2340.150 2.680 ;
        RECT 2341.270 2.310 2356.710 2.680 ;
        RECT 2357.830 2.310 2374.190 2.680 ;
        RECT 2375.310 2.310 2391.670 2.680 ;
        RECT 2392.790 2.310 2409.150 2.680 ;
        RECT 2410.270 2.310 2426.630 2.680 ;
        RECT 2427.750 2.310 2444.110 2.680 ;
        RECT 2445.230 2.310 2461.590 2.680 ;
        RECT 2462.710 2.310 2479.070 2.680 ;
        RECT 2480.190 2.310 2496.550 2.680 ;
        RECT 2497.670 2.310 2514.030 2.680 ;
        RECT 2515.150 2.310 2531.510 2.680 ;
        RECT 2532.630 2.310 2548.990 2.680 ;
        RECT 2550.110 2.310 2566.470 2.680 ;
        RECT 2567.590 2.310 2583.950 2.680 ;
        RECT 2585.070 2.310 2601.430 2.680 ;
        RECT 2602.550 2.310 2618.910 2.680 ;
        RECT 2620.030 2.310 2636.390 2.680 ;
        RECT 2637.510 2.310 2653.870 2.680 ;
        RECT 2654.990 2.310 2671.350 2.680 ;
        RECT 2672.470 2.310 2688.830 2.680 ;
        RECT 2689.950 2.310 2706.310 2.680 ;
        RECT 2707.430 2.310 2723.790 2.680 ;
        RECT 2724.910 2.310 2741.270 2.680 ;
        RECT 2742.390 2.310 2758.750 2.680 ;
        RECT 2759.870 2.310 2776.230 2.680 ;
        RECT 2777.350 2.310 2793.710 2.680 ;
        RECT 2794.830 2.310 2811.190 2.680 ;
        RECT 2812.310 2.310 2828.670 2.680 ;
        RECT 2829.790 2.310 2846.150 2.680 ;
        RECT 2847.270 2.310 2863.630 2.680 ;
        RECT 2864.750 2.310 2881.110 2.680 ;
        RECT 2882.230 2.310 2898.590 2.680 ;
        RECT 2899.710 2.310 2916.070 2.680 ;
      LAYER met3 ;
        RECT 2.800 3509.500 2917.600 3510.665 ;
        RECT 2.400 3507.420 2917.600 3509.500 ;
        RECT 2.400 3505.420 2917.200 3507.420 ;
        RECT 2.400 3485.660 2917.600 3505.420 ;
        RECT 2.800 3483.660 2917.600 3485.660 ;
        RECT 2.400 3481.580 2917.600 3483.660 ;
        RECT 2.400 3479.580 2917.200 3481.580 ;
        RECT 2.400 3461.180 2917.600 3479.580 ;
        RECT 2.800 3459.180 2917.600 3461.180 ;
        RECT 2.400 3455.740 2917.600 3459.180 ;
        RECT 2.400 3453.740 2917.200 3455.740 ;
        RECT 2.400 3435.340 2917.600 3453.740 ;
        RECT 2.800 3433.340 2917.600 3435.340 ;
        RECT 2.400 3429.900 2917.600 3433.340 ;
        RECT 2.400 3427.900 2917.200 3429.900 ;
        RECT 2.400 3409.500 2917.600 3427.900 ;
        RECT 2.800 3407.500 2917.600 3409.500 ;
        RECT 2.400 3404.060 2917.600 3407.500 ;
        RECT 2.400 3402.060 2917.200 3404.060 ;
        RECT 2.400 3383.660 2917.600 3402.060 ;
        RECT 2.800 3381.660 2917.600 3383.660 ;
        RECT 2.400 3378.220 2917.600 3381.660 ;
        RECT 2.400 3376.220 2917.200 3378.220 ;
        RECT 2.400 3357.820 2917.600 3376.220 ;
        RECT 2.800 3355.820 2917.600 3357.820 ;
        RECT 2.400 3352.380 2917.600 3355.820 ;
        RECT 2.400 3350.380 2917.200 3352.380 ;
        RECT 2.400 3331.980 2917.600 3350.380 ;
        RECT 2.800 3329.980 2917.600 3331.980 ;
        RECT 2.400 3326.540 2917.600 3329.980 ;
        RECT 2.400 3324.540 2917.200 3326.540 ;
        RECT 2.400 3306.140 2917.600 3324.540 ;
        RECT 2.800 3304.140 2917.600 3306.140 ;
        RECT 2.400 3300.700 2917.600 3304.140 ;
        RECT 2.400 3298.700 2917.200 3300.700 ;
        RECT 2.400 3280.300 2917.600 3298.700 ;
        RECT 2.800 3278.300 2917.600 3280.300 ;
        RECT 2.400 3274.860 2917.600 3278.300 ;
        RECT 2.400 3272.860 2917.200 3274.860 ;
        RECT 2.400 3254.460 2917.600 3272.860 ;
        RECT 2.800 3252.460 2917.600 3254.460 ;
        RECT 2.400 3249.020 2917.600 3252.460 ;
        RECT 2.400 3247.020 2917.200 3249.020 ;
        RECT 2.400 3228.620 2917.600 3247.020 ;
        RECT 2.800 3226.620 2917.600 3228.620 ;
        RECT 2.400 3223.180 2917.600 3226.620 ;
        RECT 2.400 3221.180 2917.200 3223.180 ;
        RECT 2.400 3202.780 2917.600 3221.180 ;
        RECT 2.800 3200.780 2917.600 3202.780 ;
        RECT 2.400 3197.340 2917.600 3200.780 ;
        RECT 2.400 3195.340 2917.200 3197.340 ;
        RECT 2.400 3176.940 2917.600 3195.340 ;
        RECT 2.800 3174.940 2917.600 3176.940 ;
        RECT 2.400 3171.500 2917.600 3174.940 ;
        RECT 2.400 3169.500 2917.200 3171.500 ;
        RECT 2.400 3151.100 2917.600 3169.500 ;
        RECT 2.800 3149.100 2917.600 3151.100 ;
        RECT 2.400 3145.660 2917.600 3149.100 ;
        RECT 2.400 3143.660 2917.200 3145.660 ;
        RECT 2.400 3125.260 2917.600 3143.660 ;
        RECT 2.800 3123.260 2917.600 3125.260 ;
        RECT 2.400 3119.820 2917.600 3123.260 ;
        RECT 2.400 3117.820 2917.200 3119.820 ;
        RECT 2.400 3099.420 2917.600 3117.820 ;
        RECT 2.800 3097.420 2917.600 3099.420 ;
        RECT 2.400 3093.980 2917.600 3097.420 ;
        RECT 2.400 3091.980 2917.200 3093.980 ;
        RECT 2.400 3073.580 2917.600 3091.980 ;
        RECT 2.800 3071.580 2917.600 3073.580 ;
        RECT 2.400 3068.140 2917.600 3071.580 ;
        RECT 2.400 3066.140 2917.200 3068.140 ;
        RECT 2.400 3047.740 2917.600 3066.140 ;
        RECT 2.800 3045.740 2917.600 3047.740 ;
        RECT 2.400 3042.300 2917.600 3045.740 ;
        RECT 2.400 3040.300 2917.200 3042.300 ;
        RECT 2.400 3021.900 2917.600 3040.300 ;
        RECT 2.800 3019.900 2917.600 3021.900 ;
        RECT 2.400 3016.460 2917.600 3019.900 ;
        RECT 2.400 3014.460 2917.200 3016.460 ;
        RECT 2.400 2996.060 2917.600 3014.460 ;
        RECT 2.800 2994.060 2917.600 2996.060 ;
        RECT 2.400 2990.620 2917.600 2994.060 ;
        RECT 2.400 2988.620 2917.200 2990.620 ;
        RECT 2.400 2970.220 2917.600 2988.620 ;
        RECT 2.800 2968.220 2917.600 2970.220 ;
        RECT 2.400 2964.780 2917.600 2968.220 ;
        RECT 2.400 2962.780 2917.200 2964.780 ;
        RECT 2.400 2944.380 2917.600 2962.780 ;
        RECT 2.800 2942.380 2917.600 2944.380 ;
        RECT 2.400 2938.940 2917.600 2942.380 ;
        RECT 2.400 2936.940 2917.200 2938.940 ;
        RECT 2.400 2918.540 2917.600 2936.940 ;
        RECT 2.800 2916.540 2917.600 2918.540 ;
        RECT 2.400 2913.100 2917.600 2916.540 ;
        RECT 2.400 2911.100 2917.200 2913.100 ;
        RECT 2.400 2892.700 2917.600 2911.100 ;
        RECT 2.800 2890.700 2917.600 2892.700 ;
        RECT 2.400 2887.260 2917.600 2890.700 ;
        RECT 2.400 2885.260 2917.200 2887.260 ;
        RECT 2.400 2866.860 2917.600 2885.260 ;
        RECT 2.800 2864.860 2917.600 2866.860 ;
        RECT 2.400 2861.420 2917.600 2864.860 ;
        RECT 2.400 2859.420 2917.200 2861.420 ;
        RECT 2.400 2841.020 2917.600 2859.420 ;
        RECT 2.800 2839.020 2917.600 2841.020 ;
        RECT 2.400 2835.580 2917.600 2839.020 ;
        RECT 2.400 2833.580 2917.200 2835.580 ;
        RECT 2.400 2815.180 2917.600 2833.580 ;
        RECT 2.800 2813.180 2917.600 2815.180 ;
        RECT 2.400 2809.740 2917.600 2813.180 ;
        RECT 2.400 2807.740 2917.200 2809.740 ;
        RECT 2.400 2789.340 2917.600 2807.740 ;
        RECT 2.800 2787.340 2917.600 2789.340 ;
        RECT 2.400 2783.900 2917.600 2787.340 ;
        RECT 2.400 2781.900 2917.200 2783.900 ;
        RECT 2.400 2763.500 2917.600 2781.900 ;
        RECT 2.800 2761.500 2917.600 2763.500 ;
        RECT 2.400 2758.060 2917.600 2761.500 ;
        RECT 2.400 2756.060 2917.200 2758.060 ;
        RECT 2.400 2737.660 2917.600 2756.060 ;
        RECT 2.800 2735.660 2917.600 2737.660 ;
        RECT 2.400 2732.220 2917.600 2735.660 ;
        RECT 2.400 2730.220 2917.200 2732.220 ;
        RECT 2.400 2711.820 2917.600 2730.220 ;
        RECT 2.800 2709.820 2917.600 2711.820 ;
        RECT 2.400 2706.380 2917.600 2709.820 ;
        RECT 2.400 2704.380 2917.200 2706.380 ;
        RECT 2.400 2685.980 2917.600 2704.380 ;
        RECT 2.800 2683.980 2917.600 2685.980 ;
        RECT 2.400 2680.540 2917.600 2683.980 ;
        RECT 2.400 2678.540 2917.200 2680.540 ;
        RECT 2.400 2660.140 2917.600 2678.540 ;
        RECT 2.800 2658.140 2917.600 2660.140 ;
        RECT 2.400 2654.700 2917.600 2658.140 ;
        RECT 2.400 2652.700 2917.200 2654.700 ;
        RECT 2.400 2634.300 2917.600 2652.700 ;
        RECT 2.800 2632.300 2917.600 2634.300 ;
        RECT 2.400 2630.220 2917.600 2632.300 ;
        RECT 2.400 2628.220 2917.200 2630.220 ;
        RECT 2.400 2608.460 2917.600 2628.220 ;
        RECT 2.800 2606.460 2917.600 2608.460 ;
        RECT 2.400 2604.380 2917.600 2606.460 ;
        RECT 2.400 2602.380 2917.200 2604.380 ;
        RECT 2.400 2582.620 2917.600 2602.380 ;
        RECT 2.800 2580.620 2917.600 2582.620 ;
        RECT 2.400 2578.540 2917.600 2580.620 ;
        RECT 2.400 2576.540 2917.200 2578.540 ;
        RECT 2.400 2556.780 2917.600 2576.540 ;
        RECT 2.800 2554.780 2917.600 2556.780 ;
        RECT 2.400 2552.700 2917.600 2554.780 ;
        RECT 2.400 2550.700 2917.200 2552.700 ;
        RECT 2.400 2530.940 2917.600 2550.700 ;
        RECT 2.800 2528.940 2917.600 2530.940 ;
        RECT 2.400 2526.860 2917.600 2528.940 ;
        RECT 2.400 2524.860 2917.200 2526.860 ;
        RECT 2.400 2505.100 2917.600 2524.860 ;
        RECT 2.800 2503.100 2917.600 2505.100 ;
        RECT 2.400 2501.020 2917.600 2503.100 ;
        RECT 2.400 2499.020 2917.200 2501.020 ;
        RECT 2.400 2479.260 2917.600 2499.020 ;
        RECT 2.800 2477.260 2917.600 2479.260 ;
        RECT 2.400 2475.180 2917.600 2477.260 ;
        RECT 2.400 2473.180 2917.200 2475.180 ;
        RECT 2.400 2453.420 2917.600 2473.180 ;
        RECT 2.800 2451.420 2917.600 2453.420 ;
        RECT 2.400 2449.340 2917.600 2451.420 ;
        RECT 2.400 2447.340 2917.200 2449.340 ;
        RECT 2.400 2427.580 2917.600 2447.340 ;
        RECT 2.800 2425.580 2917.600 2427.580 ;
        RECT 2.400 2423.500 2917.600 2425.580 ;
        RECT 2.400 2421.500 2917.200 2423.500 ;
        RECT 2.400 2401.740 2917.600 2421.500 ;
        RECT 2.800 2399.740 2917.600 2401.740 ;
        RECT 2.400 2397.660 2917.600 2399.740 ;
        RECT 2.400 2395.660 2917.200 2397.660 ;
        RECT 2.400 2375.900 2917.600 2395.660 ;
        RECT 2.800 2373.900 2917.600 2375.900 ;
        RECT 2.400 2371.820 2917.600 2373.900 ;
        RECT 2.400 2369.820 2917.200 2371.820 ;
        RECT 2.400 2350.060 2917.600 2369.820 ;
        RECT 2.800 2348.060 2917.600 2350.060 ;
        RECT 2.400 2345.980 2917.600 2348.060 ;
        RECT 2.400 2343.980 2917.200 2345.980 ;
        RECT 2.400 2324.220 2917.600 2343.980 ;
        RECT 2.800 2322.220 2917.600 2324.220 ;
        RECT 2.400 2320.140 2917.600 2322.220 ;
        RECT 2.400 2318.140 2917.200 2320.140 ;
        RECT 2.400 2298.380 2917.600 2318.140 ;
        RECT 2.800 2296.380 2917.600 2298.380 ;
        RECT 2.400 2294.300 2917.600 2296.380 ;
        RECT 2.400 2292.300 2917.200 2294.300 ;
        RECT 2.400 2272.540 2917.600 2292.300 ;
        RECT 2.800 2270.540 2917.600 2272.540 ;
        RECT 2.400 2268.460 2917.600 2270.540 ;
        RECT 2.400 2266.460 2917.200 2268.460 ;
        RECT 2.400 2246.700 2917.600 2266.460 ;
        RECT 2.800 2244.700 2917.600 2246.700 ;
        RECT 2.400 2242.620 2917.600 2244.700 ;
        RECT 2.400 2240.620 2917.200 2242.620 ;
        RECT 2.400 2220.860 2917.600 2240.620 ;
        RECT 2.800 2218.860 2917.600 2220.860 ;
        RECT 2.400 2216.780 2917.600 2218.860 ;
        RECT 2.400 2214.780 2917.200 2216.780 ;
        RECT 2.400 2195.020 2917.600 2214.780 ;
        RECT 2.800 2193.020 2917.600 2195.020 ;
        RECT 2.400 2190.940 2917.600 2193.020 ;
        RECT 2.400 2188.940 2917.200 2190.940 ;
        RECT 2.400 2169.180 2917.600 2188.940 ;
        RECT 2.800 2167.180 2917.600 2169.180 ;
        RECT 2.400 2165.100 2917.600 2167.180 ;
        RECT 2.400 2163.100 2917.200 2165.100 ;
        RECT 2.400 2143.340 2917.600 2163.100 ;
        RECT 2.800 2141.340 2917.600 2143.340 ;
        RECT 2.400 2139.260 2917.600 2141.340 ;
        RECT 2.400 2137.260 2917.200 2139.260 ;
        RECT 2.400 2117.500 2917.600 2137.260 ;
        RECT 2.800 2115.500 2917.600 2117.500 ;
        RECT 2.400 2113.420 2917.600 2115.500 ;
        RECT 2.400 2111.420 2917.200 2113.420 ;
        RECT 2.400 2091.660 2917.600 2111.420 ;
        RECT 2.800 2089.660 2917.600 2091.660 ;
        RECT 2.400 2087.580 2917.600 2089.660 ;
        RECT 2.400 2085.580 2917.200 2087.580 ;
        RECT 2.400 2065.820 2917.600 2085.580 ;
        RECT 2.800 2063.820 2917.600 2065.820 ;
        RECT 2.400 2061.740 2917.600 2063.820 ;
        RECT 2.400 2059.740 2917.200 2061.740 ;
        RECT 2.400 2039.980 2917.600 2059.740 ;
        RECT 2.800 2037.980 2917.600 2039.980 ;
        RECT 2.400 2035.900 2917.600 2037.980 ;
        RECT 2.400 2033.900 2917.200 2035.900 ;
        RECT 2.400 2014.140 2917.600 2033.900 ;
        RECT 2.800 2012.140 2917.600 2014.140 ;
        RECT 2.400 2010.060 2917.600 2012.140 ;
        RECT 2.400 2008.060 2917.200 2010.060 ;
        RECT 2.400 1988.300 2917.600 2008.060 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1984.220 2917.600 1986.300 ;
        RECT 2.400 1982.220 2917.200 1984.220 ;
        RECT 2.400 1962.460 2917.600 1982.220 ;
        RECT 2.800 1960.460 2917.600 1962.460 ;
        RECT 2.400 1958.380 2917.600 1960.460 ;
        RECT 2.400 1956.380 2917.200 1958.380 ;
        RECT 2.400 1936.620 2917.600 1956.380 ;
        RECT 2.800 1934.620 2917.600 1936.620 ;
        RECT 2.400 1932.540 2917.600 1934.620 ;
        RECT 2.400 1930.540 2917.200 1932.540 ;
        RECT 2.400 1910.780 2917.600 1930.540 ;
        RECT 2.800 1908.780 2917.600 1910.780 ;
        RECT 2.400 1906.700 2917.600 1908.780 ;
        RECT 2.400 1904.700 2917.200 1906.700 ;
        RECT 2.400 1884.940 2917.600 1904.700 ;
        RECT 2.800 1882.940 2917.600 1884.940 ;
        RECT 2.400 1880.860 2917.600 1882.940 ;
        RECT 2.400 1878.860 2917.200 1880.860 ;
        RECT 2.400 1859.100 2917.600 1878.860 ;
        RECT 2.800 1857.100 2917.600 1859.100 ;
        RECT 2.400 1855.020 2917.600 1857.100 ;
        RECT 2.400 1853.020 2917.200 1855.020 ;
        RECT 2.400 1833.260 2917.600 1853.020 ;
        RECT 2.800 1831.260 2917.600 1833.260 ;
        RECT 2.400 1829.180 2917.600 1831.260 ;
        RECT 2.400 1827.180 2917.200 1829.180 ;
        RECT 2.400 1807.420 2917.600 1827.180 ;
        RECT 2.800 1805.420 2917.600 1807.420 ;
        RECT 2.400 1803.340 2917.600 1805.420 ;
        RECT 2.400 1801.340 2917.200 1803.340 ;
        RECT 2.400 1781.580 2917.600 1801.340 ;
        RECT 2.800 1779.580 2917.600 1781.580 ;
        RECT 2.400 1777.500 2917.600 1779.580 ;
        RECT 2.400 1775.500 2917.200 1777.500 ;
        RECT 2.400 1755.740 2917.600 1775.500 ;
        RECT 2.800 1753.740 2917.600 1755.740 ;
        RECT 2.400 1751.660 2917.600 1753.740 ;
        RECT 2.400 1749.660 2917.200 1751.660 ;
        RECT 2.400 1731.260 2917.600 1749.660 ;
        RECT 2.800 1729.260 2917.600 1731.260 ;
        RECT 2.400 1725.820 2917.600 1729.260 ;
        RECT 2.400 1723.820 2917.200 1725.820 ;
        RECT 2.400 1705.420 2917.600 1723.820 ;
        RECT 2.800 1703.420 2917.600 1705.420 ;
        RECT 2.400 1699.980 2917.600 1703.420 ;
        RECT 2.400 1697.980 2917.200 1699.980 ;
        RECT 2.400 1679.580 2917.600 1697.980 ;
        RECT 2.800 1677.580 2917.600 1679.580 ;
        RECT 2.400 1674.140 2917.600 1677.580 ;
        RECT 2.400 1672.140 2917.200 1674.140 ;
        RECT 2.400 1653.740 2917.600 1672.140 ;
        RECT 2.800 1651.740 2917.600 1653.740 ;
        RECT 2.400 1648.300 2917.600 1651.740 ;
        RECT 2.400 1646.300 2917.200 1648.300 ;
        RECT 2.400 1627.900 2917.600 1646.300 ;
        RECT 2.800 1625.900 2917.600 1627.900 ;
        RECT 2.400 1622.460 2917.600 1625.900 ;
        RECT 2.400 1620.460 2917.200 1622.460 ;
        RECT 2.400 1602.060 2917.600 1620.460 ;
        RECT 2.800 1600.060 2917.600 1602.060 ;
        RECT 2.400 1596.620 2917.600 1600.060 ;
        RECT 2.400 1594.620 2917.200 1596.620 ;
        RECT 2.400 1576.220 2917.600 1594.620 ;
        RECT 2.800 1574.220 2917.600 1576.220 ;
        RECT 2.400 1570.780 2917.600 1574.220 ;
        RECT 2.400 1568.780 2917.200 1570.780 ;
        RECT 2.400 1550.380 2917.600 1568.780 ;
        RECT 2.800 1548.380 2917.600 1550.380 ;
        RECT 2.400 1544.940 2917.600 1548.380 ;
        RECT 2.400 1542.940 2917.200 1544.940 ;
        RECT 2.400 1524.540 2917.600 1542.940 ;
        RECT 2.800 1522.540 2917.600 1524.540 ;
        RECT 2.400 1519.100 2917.600 1522.540 ;
        RECT 2.400 1517.100 2917.200 1519.100 ;
        RECT 2.400 1498.700 2917.600 1517.100 ;
        RECT 2.800 1496.700 2917.600 1498.700 ;
        RECT 2.400 1493.260 2917.600 1496.700 ;
        RECT 2.400 1491.260 2917.200 1493.260 ;
        RECT 2.400 1472.860 2917.600 1491.260 ;
        RECT 2.800 1470.860 2917.600 1472.860 ;
        RECT 2.400 1467.420 2917.600 1470.860 ;
        RECT 2.400 1465.420 2917.200 1467.420 ;
        RECT 2.400 1447.020 2917.600 1465.420 ;
        RECT 2.800 1445.020 2917.600 1447.020 ;
        RECT 2.400 1441.580 2917.600 1445.020 ;
        RECT 2.400 1439.580 2917.200 1441.580 ;
        RECT 2.400 1421.180 2917.600 1439.580 ;
        RECT 2.800 1419.180 2917.600 1421.180 ;
        RECT 2.400 1415.740 2917.600 1419.180 ;
        RECT 2.400 1413.740 2917.200 1415.740 ;
        RECT 2.400 1395.340 2917.600 1413.740 ;
        RECT 2.800 1393.340 2917.600 1395.340 ;
        RECT 2.400 1389.900 2917.600 1393.340 ;
        RECT 2.400 1387.900 2917.200 1389.900 ;
        RECT 2.400 1369.500 2917.600 1387.900 ;
        RECT 2.800 1367.500 2917.600 1369.500 ;
        RECT 2.400 1364.060 2917.600 1367.500 ;
        RECT 2.400 1362.060 2917.200 1364.060 ;
        RECT 2.400 1343.660 2917.600 1362.060 ;
        RECT 2.800 1341.660 2917.600 1343.660 ;
        RECT 2.400 1338.220 2917.600 1341.660 ;
        RECT 2.400 1336.220 2917.200 1338.220 ;
        RECT 2.400 1317.820 2917.600 1336.220 ;
        RECT 2.800 1315.820 2917.600 1317.820 ;
        RECT 2.400 1312.380 2917.600 1315.820 ;
        RECT 2.400 1310.380 2917.200 1312.380 ;
        RECT 2.400 1291.980 2917.600 1310.380 ;
        RECT 2.800 1289.980 2917.600 1291.980 ;
        RECT 2.400 1286.540 2917.600 1289.980 ;
        RECT 2.400 1284.540 2917.200 1286.540 ;
        RECT 2.400 1266.140 2917.600 1284.540 ;
        RECT 2.800 1264.140 2917.600 1266.140 ;
        RECT 2.400 1260.700 2917.600 1264.140 ;
        RECT 2.400 1258.700 2917.200 1260.700 ;
        RECT 2.400 1240.300 2917.600 1258.700 ;
        RECT 2.800 1238.300 2917.600 1240.300 ;
        RECT 2.400 1234.860 2917.600 1238.300 ;
        RECT 2.400 1232.860 2917.200 1234.860 ;
        RECT 2.400 1214.460 2917.600 1232.860 ;
        RECT 2.800 1212.460 2917.600 1214.460 ;
        RECT 2.400 1209.020 2917.600 1212.460 ;
        RECT 2.400 1207.020 2917.200 1209.020 ;
        RECT 2.400 1188.620 2917.600 1207.020 ;
        RECT 2.800 1186.620 2917.600 1188.620 ;
        RECT 2.400 1183.180 2917.600 1186.620 ;
        RECT 2.400 1181.180 2917.200 1183.180 ;
        RECT 2.400 1162.780 2917.600 1181.180 ;
        RECT 2.800 1160.780 2917.600 1162.780 ;
        RECT 2.400 1157.340 2917.600 1160.780 ;
        RECT 2.400 1155.340 2917.200 1157.340 ;
        RECT 2.400 1136.940 2917.600 1155.340 ;
        RECT 2.800 1134.940 2917.600 1136.940 ;
        RECT 2.400 1131.500 2917.600 1134.940 ;
        RECT 2.400 1129.500 2917.200 1131.500 ;
        RECT 2.400 1111.100 2917.600 1129.500 ;
        RECT 2.800 1109.100 2917.600 1111.100 ;
        RECT 2.400 1105.660 2917.600 1109.100 ;
        RECT 2.400 1103.660 2917.200 1105.660 ;
        RECT 2.400 1085.260 2917.600 1103.660 ;
        RECT 2.800 1083.260 2917.600 1085.260 ;
        RECT 2.400 1079.820 2917.600 1083.260 ;
        RECT 2.400 1077.820 2917.200 1079.820 ;
        RECT 2.400 1059.420 2917.600 1077.820 ;
        RECT 2.800 1057.420 2917.600 1059.420 ;
        RECT 2.400 1053.980 2917.600 1057.420 ;
        RECT 2.400 1051.980 2917.200 1053.980 ;
        RECT 2.400 1033.580 2917.600 1051.980 ;
        RECT 2.800 1031.580 2917.600 1033.580 ;
        RECT 2.400 1028.140 2917.600 1031.580 ;
        RECT 2.400 1026.140 2917.200 1028.140 ;
        RECT 2.400 1007.740 2917.600 1026.140 ;
        RECT 2.800 1005.740 2917.600 1007.740 ;
        RECT 2.400 1002.300 2917.600 1005.740 ;
        RECT 2.400 1000.300 2917.200 1002.300 ;
        RECT 2.400 981.900 2917.600 1000.300 ;
        RECT 2.800 979.900 2917.600 981.900 ;
        RECT 2.400 976.460 2917.600 979.900 ;
        RECT 2.400 974.460 2917.200 976.460 ;
        RECT 2.400 956.060 2917.600 974.460 ;
        RECT 2.800 954.060 2917.600 956.060 ;
        RECT 2.400 950.620 2917.600 954.060 ;
        RECT 2.400 948.620 2917.200 950.620 ;
        RECT 2.400 930.220 2917.600 948.620 ;
        RECT 2.800 928.220 2917.600 930.220 ;
        RECT 2.400 924.780 2917.600 928.220 ;
        RECT 2.400 922.780 2917.200 924.780 ;
        RECT 2.400 904.380 2917.600 922.780 ;
        RECT 2.800 902.380 2917.600 904.380 ;
        RECT 2.400 900.300 2917.600 902.380 ;
        RECT 2.400 898.300 2917.200 900.300 ;
        RECT 2.400 878.540 2917.600 898.300 ;
        RECT 2.800 876.540 2917.600 878.540 ;
        RECT 2.400 874.460 2917.600 876.540 ;
        RECT 2.400 872.460 2917.200 874.460 ;
        RECT 2.400 852.700 2917.600 872.460 ;
        RECT 2.800 850.700 2917.600 852.700 ;
        RECT 2.400 848.620 2917.600 850.700 ;
        RECT 2.400 846.620 2917.200 848.620 ;
        RECT 2.400 826.860 2917.600 846.620 ;
        RECT 2.800 824.860 2917.600 826.860 ;
        RECT 2.400 822.780 2917.600 824.860 ;
        RECT 2.400 820.780 2917.200 822.780 ;
        RECT 2.400 801.020 2917.600 820.780 ;
        RECT 2.800 799.020 2917.600 801.020 ;
        RECT 2.400 796.940 2917.600 799.020 ;
        RECT 2.400 794.940 2917.200 796.940 ;
        RECT 2.400 775.180 2917.600 794.940 ;
        RECT 2.800 773.180 2917.600 775.180 ;
        RECT 2.400 771.100 2917.600 773.180 ;
        RECT 2.400 769.100 2917.200 771.100 ;
        RECT 2.400 749.340 2917.600 769.100 ;
        RECT 2.800 747.340 2917.600 749.340 ;
        RECT 2.400 745.260 2917.600 747.340 ;
        RECT 2.400 743.260 2917.200 745.260 ;
        RECT 2.400 723.500 2917.600 743.260 ;
        RECT 2.800 721.500 2917.600 723.500 ;
        RECT 2.400 719.420 2917.600 721.500 ;
        RECT 2.400 717.420 2917.200 719.420 ;
        RECT 2.400 697.660 2917.600 717.420 ;
        RECT 2.800 695.660 2917.600 697.660 ;
        RECT 2.400 693.580 2917.600 695.660 ;
        RECT 2.400 691.580 2917.200 693.580 ;
        RECT 2.400 671.820 2917.600 691.580 ;
        RECT 2.800 669.820 2917.600 671.820 ;
        RECT 2.400 667.740 2917.600 669.820 ;
        RECT 2.400 665.740 2917.200 667.740 ;
        RECT 2.400 645.980 2917.600 665.740 ;
        RECT 2.800 643.980 2917.600 645.980 ;
        RECT 2.400 641.900 2917.600 643.980 ;
        RECT 2.400 639.900 2917.200 641.900 ;
        RECT 2.400 620.140 2917.600 639.900 ;
        RECT 2.800 618.140 2917.600 620.140 ;
        RECT 2.400 616.060 2917.600 618.140 ;
        RECT 2.400 614.060 2917.200 616.060 ;
        RECT 2.400 594.300 2917.600 614.060 ;
        RECT 2.800 592.300 2917.600 594.300 ;
        RECT 2.400 590.220 2917.600 592.300 ;
        RECT 2.400 588.220 2917.200 590.220 ;
        RECT 2.400 568.460 2917.600 588.220 ;
        RECT 2.800 566.460 2917.600 568.460 ;
        RECT 2.400 564.380 2917.600 566.460 ;
        RECT 2.400 562.380 2917.200 564.380 ;
        RECT 2.400 542.620 2917.600 562.380 ;
        RECT 2.800 540.620 2917.600 542.620 ;
        RECT 2.400 538.540 2917.600 540.620 ;
        RECT 2.400 536.540 2917.200 538.540 ;
        RECT 2.400 516.780 2917.600 536.540 ;
        RECT 2.800 514.780 2917.600 516.780 ;
        RECT 2.400 512.700 2917.600 514.780 ;
        RECT 2.400 510.700 2917.200 512.700 ;
        RECT 2.400 490.940 2917.600 510.700 ;
        RECT 2.800 488.940 2917.600 490.940 ;
        RECT 2.400 486.860 2917.600 488.940 ;
        RECT 2.400 484.860 2917.200 486.860 ;
        RECT 2.400 465.100 2917.600 484.860 ;
        RECT 2.800 463.100 2917.600 465.100 ;
        RECT 2.400 461.020 2917.600 463.100 ;
        RECT 2.400 459.020 2917.200 461.020 ;
        RECT 2.400 439.260 2917.600 459.020 ;
        RECT 2.800 437.260 2917.600 439.260 ;
        RECT 2.400 435.180 2917.600 437.260 ;
        RECT 2.400 433.180 2917.200 435.180 ;
        RECT 2.400 413.420 2917.600 433.180 ;
        RECT 2.800 411.420 2917.600 413.420 ;
        RECT 2.400 409.340 2917.600 411.420 ;
        RECT 2.400 407.340 2917.200 409.340 ;
        RECT 2.400 387.580 2917.600 407.340 ;
        RECT 2.800 385.580 2917.600 387.580 ;
        RECT 2.400 383.500 2917.600 385.580 ;
        RECT 2.400 381.500 2917.200 383.500 ;
        RECT 2.400 361.740 2917.600 381.500 ;
        RECT 2.800 359.740 2917.600 361.740 ;
        RECT 2.400 357.660 2917.600 359.740 ;
        RECT 2.400 355.660 2917.200 357.660 ;
        RECT 2.400 335.900 2917.600 355.660 ;
        RECT 2.800 333.900 2917.600 335.900 ;
        RECT 2.400 331.820 2917.600 333.900 ;
        RECT 2.400 329.820 2917.200 331.820 ;
        RECT 2.400 310.060 2917.600 329.820 ;
        RECT 2.800 308.060 2917.600 310.060 ;
        RECT 2.400 305.980 2917.600 308.060 ;
        RECT 2.400 303.980 2917.200 305.980 ;
        RECT 2.400 284.220 2917.600 303.980 ;
        RECT 2.800 282.220 2917.600 284.220 ;
        RECT 2.400 280.140 2917.600 282.220 ;
        RECT 2.400 278.140 2917.200 280.140 ;
        RECT 2.400 258.380 2917.600 278.140 ;
        RECT 2.800 256.380 2917.600 258.380 ;
        RECT 2.400 254.300 2917.600 256.380 ;
        RECT 2.400 252.300 2917.200 254.300 ;
        RECT 2.400 232.540 2917.600 252.300 ;
        RECT 2.800 230.540 2917.600 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.400 226.460 2917.200 228.460 ;
        RECT 2.400 206.700 2917.600 226.460 ;
        RECT 2.800 204.700 2917.600 206.700 ;
        RECT 2.400 202.620 2917.600 204.700 ;
        RECT 2.400 200.620 2917.200 202.620 ;
        RECT 2.400 180.860 2917.600 200.620 ;
        RECT 2.800 178.860 2917.600 180.860 ;
        RECT 2.400 176.780 2917.600 178.860 ;
        RECT 2.400 174.780 2917.200 176.780 ;
        RECT 2.400 155.020 2917.600 174.780 ;
        RECT 2.800 153.020 2917.600 155.020 ;
        RECT 2.400 150.940 2917.600 153.020 ;
        RECT 2.400 148.940 2917.200 150.940 ;
        RECT 2.400 129.180 2917.600 148.940 ;
        RECT 2.800 127.180 2917.600 129.180 ;
        RECT 2.400 125.100 2917.600 127.180 ;
        RECT 2.400 123.100 2917.200 125.100 ;
        RECT 2.400 103.340 2917.600 123.100 ;
        RECT 2.800 101.340 2917.600 103.340 ;
        RECT 2.400 99.260 2917.600 101.340 ;
        RECT 2.400 97.260 2917.200 99.260 ;
        RECT 2.400 77.500 2917.600 97.260 ;
        RECT 2.800 75.500 2917.600 77.500 ;
        RECT 2.400 73.420 2917.600 75.500 ;
        RECT 2.400 71.420 2917.200 73.420 ;
        RECT 2.400 51.660 2917.600 71.420 ;
        RECT 2.800 49.660 2917.600 51.660 ;
        RECT 2.400 47.580 2917.600 49.660 ;
        RECT 2.400 45.580 2917.200 47.580 ;
        RECT 2.400 25.820 2917.600 45.580 ;
        RECT 2.800 23.820 2917.600 25.820 ;
        RECT 2.400 21.740 2917.600 23.820 ;
        RECT 2.400 19.740 2917.200 21.740 ;
        RECT 2.400 15.135 2917.600 19.740 ;
      LAYER met4 ;
        RECT 521.040 15.135 1981.840 3504.545 ;
  END
END top
END LIBRARY

