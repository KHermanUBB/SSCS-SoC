magic
tech sky130A
magscale 1 2
timestamp 1633795376
<< locali >>
rect 284217 610283 284251 610589
rect 50997 599131 51031 599233
rect 80989 565879 81023 566049
rect 16129 561527 16163 561629
rect 12357 524603 12391 525045
rect 350917 524739 350951 525045
rect 248521 506923 248555 507365
rect 250269 506787 250303 507161
rect 256065 496043 256099 496349
rect 278697 491623 278731 492133
rect 432429 469727 432463 469829
rect 112637 467143 112671 467449
rect 154037 443139 154071 443581
rect 42165 439467 42199 439773
rect 44005 439331 44039 439705
rect 332057 423147 332091 423521
rect 28365 422807 28399 422909
rect 32045 422807 32079 423045
rect 279709 415395 279743 415429
rect 279709 415361 279893 415395
rect 57805 409275 57839 409513
rect 23397 394723 23431 394825
rect 198013 383911 198047 384149
rect 199393 383639 199427 384761
rect 200589 383911 200623 384149
rect 200405 383639 200439 383809
rect 143457 365347 143491 365449
rect 5365 348483 5399 348585
rect 311725 333999 311759 334305
rect 314485 334305 314795 334339
rect 314485 334203 314519 334305
rect 314761 334271 314795 334305
rect 314669 334067 314703 334237
rect 251189 329035 251223 329341
rect 426449 308567 426483 308669
rect 49893 304351 49927 304861
rect 112821 295647 112855 295817
rect 375297 270691 375331 271065
rect 126069 260899 126103 261001
rect 265725 223363 265759 223533
rect 260849 223159 260883 223261
rect 75837 220439 75871 220609
rect 78965 220439 78999 220541
rect 96169 220439 96203 220541
rect 97181 220439 97215 220541
rect 124137 219895 124171 220609
rect 9505 217719 9539 219045
rect 11805 218467 11839 219521
rect 12817 218535 12851 219521
rect 16221 218603 16255 219521
rect 17233 218671 17267 219521
rect 22937 218807 22971 219317
rect 53757 218807 53791 219453
rect 78137 218875 78171 219317
rect 96077 218875 96111 219521
rect 114385 218263 114419 219317
rect 128369 219011 128403 220609
rect 128461 218943 128495 220677
rect 129105 219963 129139 220541
rect 133797 220167 133831 220609
rect 167101 220031 167135 220609
rect 178049 220099 178083 220405
rect 204821 219895 204855 220473
rect 257997 219963 258031 220609
rect 258089 220099 258123 220405
rect 266645 219895 266679 220677
rect 267013 220099 267047 220609
rect 272441 220099 272475 220541
rect 272533 220371 272567 220541
rect 254961 219691 254995 219793
rect 266737 219691 266771 219861
rect 287621 219487 287655 220609
rect 232973 218739 233007 219317
rect 248337 218739 248371 219317
rect 370881 216767 370915 216869
rect 370973 216835 371007 216937
rect 322489 152167 322523 152405
rect 322339 152133 322523 152167
rect 9597 142171 9631 145129
rect 9781 136391 9815 142273
rect 7481 135371 7515 136357
rect 248889 120683 248923 120785
rect 299673 120683 299707 120853
rect 239229 119969 239447 120003
rect 239229 119935 239263 119969
rect 35725 119051 35759 119425
rect 75745 119323 75779 119765
rect 80989 119323 81023 119833
rect 145297 118711 145331 119425
rect 156613 119391 156647 119901
rect 166273 119391 166307 119901
rect 233893 119663 233927 119901
rect 239321 119459 239355 119901
rect 239229 119425 239355 119459
rect 233893 119391 233927 119425
rect 239229 119391 239263 119425
rect 233893 119357 234077 119391
rect 239413 119391 239447 119969
rect 239413 119357 239505 119391
rect 214481 118983 214515 119357
rect 216321 118983 216355 119289
rect 233341 119255 233375 119357
rect 238309 118779 238343 119289
rect 239597 119187 239631 120037
rect 248521 119391 248555 119629
rect 248463 119357 248555 119391
rect 253121 119323 253155 119493
rect 239321 118847 239355 119153
rect 248521 118847 248555 119017
rect 253949 118847 253983 119153
rect 253949 118813 254225 118847
rect 254501 118779 254535 119085
rect 255237 118915 255271 119425
rect 258641 119323 258675 119697
rect 258733 119255 258767 119425
rect 289829 119391 289863 119969
rect 289921 119663 289955 119969
rect 290013 119765 290783 119799
rect 290013 119731 290047 119765
rect 290749 119731 290783 119765
rect 291853 119663 291887 119969
rect 291945 119527 291979 119969
rect 307711 119765 308263 119799
rect 308229 119731 308263 119765
rect 301605 119119 301639 119289
rect 253983 118745 254535 118779
rect 258917 118779 258951 119085
rect 289311 118813 289461 118847
rect 291853 118779 291887 118881
rect 291945 118779 291979 119085
rect 297925 118915 297959 119085
rect 307677 118847 307711 119289
rect 308229 119051 308263 119085
rect 307861 119017 308263 119051
rect 307861 118779 307895 119017
rect 307527 118745 307895 118779
rect 28641 110755 28675 111129
rect 50997 110619 51031 110721
rect 82829 110687 82863 110857
rect 84025 110687 84059 111401
rect 106289 110687 106323 111061
rect 108313 110687 108347 111061
rect 108405 110551 108439 111061
rect 132049 110551 132083 111741
rect 166273 110755 166307 111469
rect 170505 110755 170539 111469
rect 173817 111367 173851 111469
rect 173909 111095 173943 111333
rect 178969 111231 179003 111469
rect 179061 111367 179095 111673
rect 179153 111163 179187 111333
rect 179613 111163 179647 111197
rect 179613 111129 179981 111163
rect 170413 110551 170447 110721
rect 178601 110211 178635 110721
rect 178693 110279 178727 110789
rect 181085 110279 181119 110789
rect 183109 110755 183143 111197
rect 183385 111095 183419 111673
rect 183201 110211 183235 110721
rect 183293 110687 183327 111061
rect 187801 110959 187835 111469
rect 191021 111231 191055 111333
rect 190101 110891 190135 111197
rect 190929 111163 190963 111197
rect 190929 111129 191055 111163
rect 191021 110619 191055 111129
rect 194885 110891 194919 111469
rect 202521 110483 202555 111333
rect 212641 110823 212675 111197
rect 221657 110755 221691 111537
rect 221657 110721 221749 110755
rect 221657 110279 221691 110653
rect 222761 110619 222795 111401
rect 326813 111231 326847 111741
rect 222945 110823 222979 111197
rect 272441 110959 272475 111129
rect 274097 110959 274131 111129
rect 274189 110687 274223 111129
rect 327917 111095 327951 111741
rect 328009 111231 328043 111741
rect 329757 111231 329791 111809
rect 224969 110483 225003 110653
rect 282101 110687 282135 110925
rect 286425 110687 286459 110925
rect 225245 110279 225279 110653
rect 286517 110483 286551 110653
rect 380909 85663 380943 85765
rect 340613 45951 340647 46053
rect 392501 34527 392535 35037
rect 478797 13719 478831 13821
rect 35725 9163 35759 9537
rect 66177 8347 66211 9537
rect 76757 8551 76791 9401
rect 77493 8619 77527 9537
rect 115857 9367 115891 9537
rect 115949 8959 115983 9333
rect 116041 8823 116075 9469
rect 121469 9367 121503 9469
rect 120089 8755 120123 9333
rect 138397 9027 138431 9469
rect 142169 9299 142203 9401
rect 148517 8415 148551 9333
rect 148977 8755 149011 9469
rect 150357 8891 150391 9061
rect 150449 8687 150483 9333
rect 150541 9095 150575 9469
rect 151737 9367 151771 9537
rect 152933 8687 152967 9537
rect 153025 8891 153059 9469
rect 161489 9231 161523 9333
rect 154037 9095 154071 9197
rect 153117 8415 153151 8857
rect 168389 8619 168423 9333
rect 168481 9095 168515 9197
rect 170321 9095 170355 9333
rect 185409 9299 185443 9673
rect 185501 9367 185535 9537
rect 186237 9299 186271 9673
rect 191205 9367 191239 9537
rect 233893 9231 233927 9401
rect 168297 8415 168331 8585
rect 170321 8415 170355 9061
rect 171793 8619 171827 9197
rect 233801 8823 233835 9061
rect 241529 8891 241563 9537
rect 243461 8891 243495 9401
rect 230397 8619 230431 8789
rect 245117 8483 245151 9401
rect 245577 8483 245611 9537
rect 247877 8415 247911 9537
rect 266829 9435 266863 9469
rect 266829 9401 267105 9435
rect 258641 9367 258675 9401
rect 258641 9333 258917 9367
rect 253121 8823 253155 9061
rect 253305 8891 253339 9197
rect 263643 9129 263827 9163
rect 253213 8619 253247 8789
rect 253397 8483 253431 8857
rect 258641 8823 258675 9061
rect 261677 9061 261769 9095
rect 261677 8823 261711 9061
rect 258549 8619 258583 8789
rect 261769 8619 261803 8789
rect 263701 8619 263735 9061
rect 263793 8551 263827 9129
rect 267197 8755 267231 9333
rect 268393 8619 268427 8789
rect 271429 8551 271463 9469
rect 263643 8449 263885 8483
rect 271521 8415 271555 9673
rect 277501 9469 277593 9503
rect 273729 8619 273763 9333
rect 277501 9095 277535 9469
rect 277443 9061 277535 9095
rect 277777 8415 277811 8585
rect 278053 8415 278087 9673
rect 278145 9299 278179 9877
rect 280813 9095 280847 9265
rect 282193 9231 282227 9469
rect 282101 9163 282135 9197
rect 282285 9163 282319 9469
rect 282101 9129 282319 9163
rect 280813 9061 280997 9095
rect 279341 8755 279375 8789
rect 279191 8721 279375 8755
rect 282193 8755 282227 9061
rect 282285 8687 282319 8721
rect 282101 8653 282319 8687
rect 282101 8415 282135 8653
rect 282193 8415 282227 8517
rect 310989 3383 311023 4029
rect 318717 3383 318751 4029
rect 312093 3043 312127 3349
rect 498209 3247 498243 45917
<< viali >>
rect 364257 614941 364291 614975
rect 167561 613921 167595 613955
rect 167285 613853 167319 613887
rect 167469 613853 167503 613887
rect 167653 613853 167687 613887
rect 167745 613853 167779 613887
rect 167929 613717 167963 613751
rect 376217 611677 376251 611711
rect 376033 611541 376067 611575
rect 283021 610589 283055 610623
rect 283169 610589 283203 610623
rect 283527 610589 283561 610623
rect 284217 610589 284251 610623
rect 283297 610521 283331 610555
rect 283389 610521 283423 610555
rect 283665 610453 283699 610487
rect 284217 610249 284251 610283
rect 200865 609501 200899 609535
rect 129657 608821 129691 608855
rect 334909 607937 334943 607971
rect 334725 607733 334759 607767
rect 200497 607325 200531 607359
rect 200405 607189 200439 607223
rect 228456 606849 228490 606883
rect 228189 606781 228223 606815
rect 229569 606645 229603 606679
rect 322213 604061 322247 604095
rect 184581 601409 184615 601443
rect 22753 600797 22787 600831
rect 23020 600729 23054 600763
rect 24133 600661 24167 600695
rect 233433 600253 233467 600287
rect 50445 599301 50479 599335
rect 50348 599233 50382 599267
rect 50537 599233 50571 599267
rect 50721 599233 50755 599267
rect 50997 599233 51031 599267
rect 50997 599097 51031 599131
rect 50169 599029 50203 599063
rect 247601 596649 247635 596683
rect 206017 596513 206051 596547
rect 205465 596309 205499 596343
rect 205833 596309 205867 596343
rect 205925 596309 205959 596343
rect 492965 591209 492999 591243
rect 494345 591005 494379 591039
rect 494078 590937 494112 590971
rect 419549 590597 419583 590631
rect 419365 590529 419399 590563
rect 419641 590325 419675 590359
rect 463433 587265 463467 587299
rect 463525 587265 463559 587299
rect 463157 587197 463191 587231
rect 463249 587061 463283 587095
rect 463709 587061 463743 587095
rect 313381 586177 313415 586211
rect 410349 585565 410383 585599
rect 106749 584681 106783 584715
rect 201601 584001 201635 584035
rect 201325 583933 201359 583967
rect 201509 583933 201543 583967
rect 201969 583797 202003 583831
rect 405933 583389 405967 583423
rect 482569 580737 482603 580771
rect 482661 580669 482695 580703
rect 482753 580669 482787 580703
rect 482201 580533 482235 580567
rect 396917 579105 396951 579139
rect 113649 579037 113683 579071
rect 396641 578969 396675 579003
rect 396273 578901 396307 578935
rect 396733 578901 396767 578935
rect 248245 578357 248279 578391
rect 423781 576929 423815 576963
rect 423413 576861 423447 576895
rect 423597 576861 423631 576895
rect 417525 576181 417559 576215
rect 196449 572033 196483 572067
rect 196716 572033 196750 572067
rect 369409 571965 369443 571999
rect 197829 571829 197863 571863
rect 236469 571081 236503 571115
rect 237582 570945 237616 570979
rect 237849 570945 237883 570979
rect 285321 570945 285355 570979
rect 376493 569245 376527 569279
rect 473737 567069 473771 567103
rect 473921 567069 473955 567103
rect 473829 566933 473863 566967
rect 78597 566185 78631 566219
rect 80989 566049 81023 566083
rect 75653 565981 75687 566015
rect 75837 565981 75871 566015
rect 75930 565959 75964 565993
rect 76022 565981 76056 566015
rect 76297 565913 76331 565947
rect 325617 565981 325651 566015
rect 325801 565981 325835 566015
rect 325525 565913 325559 565947
rect 80989 565845 81023 565879
rect 15025 561697 15059 561731
rect 15485 561697 15519 561731
rect 15209 561629 15243 561663
rect 15301 561629 15335 561663
rect 15577 561629 15611 561663
rect 16129 561629 16163 561663
rect 16129 561493 16163 561527
rect 203993 559113 204027 559147
rect 204177 558977 204211 559011
rect 204361 558909 204395 558943
rect 403449 557345 403483 557379
rect 403265 557209 403299 557243
rect 402897 557141 402931 557175
rect 403357 557141 403391 557175
rect 169953 556801 169987 556835
rect 170137 556801 170171 556835
rect 169861 556665 169895 556699
rect 304917 555101 304951 555135
rect 330861 554013 330895 554047
rect 268347 553537 268381 553571
rect 268485 553537 268519 553571
rect 268577 553537 268611 553571
rect 268760 553537 268794 553571
rect 268853 553537 268887 553571
rect 268209 553401 268243 553435
rect 434908 551837 434942 551871
rect 435280 551837 435314 551871
rect 435373 551837 435407 551871
rect 435005 551769 435039 551803
rect 435097 551769 435131 551803
rect 434729 551701 434763 551735
rect 231869 548641 231903 548675
rect 232136 548505 232170 548539
rect 233249 548437 233283 548471
rect 380633 547485 380667 547519
rect 380366 547417 380400 547451
rect 379253 547349 379287 547383
rect 121837 546805 121871 546839
rect 416605 544221 416639 544255
rect 445033 544221 445067 544255
rect 157257 543745 157291 543779
rect 157441 543745 157475 543779
rect 157625 543745 157659 543779
rect 119537 541705 119571 541739
rect 119721 541569 119755 541603
rect 119813 541569 119847 541603
rect 120089 541501 120123 541535
rect 119997 541433 120031 541467
rect 158453 540481 158487 540515
rect 158637 540481 158671 540515
rect 158729 540481 158763 540515
rect 158822 540471 158856 540505
rect 159097 540345 159131 540379
rect 59369 539393 59403 539427
rect 59461 539393 59495 539427
rect 59737 539325 59771 539359
rect 59185 539189 59219 539223
rect 59645 539189 59679 539223
rect 17325 537693 17359 537727
rect 441905 537693 441939 537727
rect 327917 536605 327951 536639
rect 331505 534633 331539 534667
rect 331321 534429 331355 534463
rect 136189 533953 136223 533987
rect 136097 533749 136131 533783
rect 342453 531573 342487 531607
rect 355609 528989 355643 529023
rect 355517 528853 355551 528887
rect 91385 528309 91419 528343
rect 13001 527901 13035 527935
rect 353953 527901 353987 527935
rect 12734 527833 12768 527867
rect 11621 527765 11655 527799
rect 376778 527425 376812 527459
rect 377045 527425 377079 527459
rect 375665 527221 375699 527255
rect 121101 526337 121135 526371
rect 121009 526133 121043 526167
rect 262781 525249 262815 525283
rect 262505 525181 262539 525215
rect 262689 525181 262723 525215
rect 351469 525181 351503 525215
rect 351745 525181 351779 525215
rect 12357 525045 12391 525079
rect 263149 525045 263183 525079
rect 350917 525045 350951 525079
rect 10885 524705 10919 524739
rect 11529 524705 11563 524739
rect 11253 524637 11287 524671
rect 11713 524637 11747 524671
rect 350917 524705 350951 524739
rect 351561 524705 351595 524739
rect 351745 524705 351779 524739
rect 12357 524569 12391 524603
rect 351469 524569 351503 524603
rect 11437 524501 11471 524535
rect 351101 524501 351135 524535
rect 291117 518721 291151 518755
rect 291209 518653 291243 518687
rect 291301 518653 291335 518687
rect 290749 518517 290783 518551
rect 319913 514845 319947 514879
rect 319821 514777 319855 514811
rect 92029 514369 92063 514403
rect 405749 514369 405783 514403
rect 405841 514301 405875 514335
rect 406025 514301 406059 514335
rect 92121 514165 92155 514199
rect 405381 514165 405415 514199
rect 46213 513961 46247 513995
rect 260665 513825 260699 513859
rect 24409 513757 24443 513791
rect 45937 513757 45971 513791
rect 46029 513757 46063 513791
rect 46213 513689 46247 513723
rect 260398 513689 260432 513723
rect 45753 513621 45787 513655
rect 259285 513621 259319 513655
rect 317337 510901 317371 510935
rect 326353 507977 326387 508011
rect 325229 507841 325263 507875
rect 426633 507841 426667 507875
rect 426817 507841 426851 507875
rect 324973 507773 325007 507807
rect 426909 507637 426943 507671
rect 247693 507433 247727 507467
rect 248521 507365 248555 507399
rect 247601 507229 247635 507263
rect 247877 507229 247911 507263
rect 247969 507229 248003 507263
rect 248153 507093 248187 507127
rect 250085 507229 250119 507263
rect 248889 507161 248923 507195
rect 250269 507161 250303 507195
rect 248521 506889 248555 506923
rect 248797 506889 248831 506923
rect 249257 506753 249291 506787
rect 250269 506753 250303 506787
rect 383945 504577 383979 504611
rect 383853 504373 383887 504407
rect 116777 502197 116811 502231
rect 420745 500769 420779 500803
rect 420929 500701 420963 500735
rect 421021 500701 421055 500735
rect 420561 500633 420595 500667
rect 420653 500633 420687 500667
rect 421205 500633 421239 500667
rect 190377 500021 190411 500055
rect 208225 498117 208259 498151
rect 208409 498117 208443 498151
rect 208593 498049 208627 498083
rect 256801 496417 256835 496451
rect 255605 496349 255639 496383
rect 256065 496349 256099 496383
rect 256341 496349 256375 496383
rect 255789 496213 255823 496247
rect 255881 496009 255915 496043
rect 256065 496009 256099 496043
rect 255697 495873 255731 495907
rect 256341 495873 256375 495907
rect 257169 495805 257203 495839
rect 204913 494581 204947 494615
rect 229109 494173 229143 494207
rect 32137 493153 32171 493187
rect 32321 493017 32355 493051
rect 32413 492949 32447 492983
rect 32781 492949 32815 492983
rect 278329 492133 278363 492167
rect 278697 492133 278731 492167
rect 276949 492065 276983 492099
rect 208501 491997 208535 492031
rect 208256 491929 208290 491963
rect 277216 491929 277250 491963
rect 207121 491861 207155 491895
rect 278697 491589 278731 491623
rect 248061 489821 248095 489855
rect 412925 489821 412959 489855
rect 248328 489753 248362 489787
rect 413170 489753 413204 489787
rect 249441 489685 249475 489719
rect 414305 489685 414339 489719
rect 470057 489141 470091 489175
rect 21465 487305 21499 487339
rect 21005 487237 21039 487271
rect 417525 487237 417559 487271
rect 21097 487169 21131 487203
rect 417800 487191 417834 487225
rect 417892 487191 417926 487225
rect 417985 487169 418019 487203
rect 418169 487169 418203 487203
rect 20913 487101 20947 487135
rect 264069 485605 264103 485639
rect 263885 485469 263919 485503
rect 263517 485333 263551 485367
rect 263701 485333 263735 485367
rect 263793 485333 263827 485367
rect 464169 484041 464203 484075
rect 464261 484041 464295 484075
rect 463985 483905 464019 483939
rect 464353 483905 464387 483939
rect 464537 483769 464571 483803
rect 382565 482409 382599 482443
rect 383945 482273 383979 482307
rect 383678 482137 383712 482171
rect 16405 480641 16439 480675
rect 16589 480573 16623 480607
rect 16221 480437 16255 480471
rect 238217 480097 238251 480131
rect 238484 479961 238518 479995
rect 239597 479893 239631 479927
rect 495357 475745 495391 475779
rect 495265 475677 495299 475711
rect 495541 475677 495575 475711
rect 495633 475677 495667 475711
rect 495817 475541 495851 475575
rect 94053 473569 94087 473603
rect 93869 473501 93903 473535
rect 202705 473501 202739 473535
rect 202889 473501 202923 473535
rect 93409 473365 93443 473399
rect 93777 473365 93811 473399
rect 203073 473365 203107 473399
rect 198657 471325 198691 471359
rect 198289 471257 198323 471291
rect 198473 471257 198507 471291
rect 149345 470849 149379 470883
rect 149612 470849 149646 470883
rect 150725 470645 150759 470679
rect 432429 469829 432463 469863
rect 432777 469761 432811 469795
rect 432429 469693 432463 469727
rect 432521 469693 432555 469727
rect 433901 469557 433935 469591
rect 112637 467449 112671 467483
rect 111901 467177 111935 467211
rect 112637 467109 112671 467143
rect 112361 467041 112395 467075
rect 194793 467041 194827 467075
rect 112085 466973 112119 467007
rect 112177 466973 112211 467007
rect 112453 466973 112487 467007
rect 195060 466905 195094 466939
rect 196173 466837 196207 466871
rect 223037 465409 223071 465443
rect 223129 465341 223163 465375
rect 223313 465341 223347 465375
rect 223865 465341 223899 465375
rect 224417 465341 224451 465375
rect 222669 465205 222703 465239
rect 362785 463709 362819 463743
rect 109785 463029 109819 463063
rect 170413 460921 170447 460955
rect 185593 457589 185627 457623
rect 254225 457181 254259 457215
rect 254133 457045 254167 457079
rect 133797 454325 133831 454359
rect 315313 453237 315347 453271
rect 53647 451265 53681 451299
rect 53757 451265 53791 451299
rect 54033 451265 54067 451299
rect 53481 451061 53515 451095
rect 53941 451061 53975 451095
rect 175933 448545 175967 448579
rect 175795 448477 175829 448511
rect 176025 448477 176059 448511
rect 175565 448409 175599 448443
rect 175657 448409 175691 448443
rect 176209 448409 176243 448443
rect 64797 447797 64831 447831
rect 112269 446913 112303 446947
rect 112361 446913 112395 446947
rect 334642 446913 334676 446947
rect 112453 446845 112487 446879
rect 334909 446845 334943 446879
rect 111901 446709 111935 446743
rect 333529 446709 333563 446743
rect 152381 443649 152415 443683
rect 423965 443649 423999 443683
rect 152473 443581 152507 443615
rect 152657 443581 152691 443615
rect 153209 443581 153243 443615
rect 153853 443581 153887 443615
rect 154037 443581 154071 443615
rect 152013 443445 152047 443479
rect 424057 443445 424091 443479
rect 152473 443105 152507 443139
rect 154037 443105 154071 443139
rect 153025 442969 153059 443003
rect 281365 442561 281399 442595
rect 376217 441949 376251 441983
rect 376125 441813 376159 441847
rect 418537 439841 418571 439875
rect 42165 439773 42199 439807
rect 42441 439773 42475 439807
rect 418445 439773 418479 439807
rect 418721 439773 418755 439807
rect 418813 439773 418847 439807
rect 43637 439705 43671 439739
rect 44005 439705 44039 439739
rect 41981 439433 42015 439467
rect 42165 439433 42199 439467
rect 43085 439433 43119 439467
rect 418997 439637 419031 439671
rect 41797 439297 41831 439331
rect 42533 439297 42567 439331
rect 44005 439297 44039 439331
rect 397101 436917 397135 436951
rect 47771 434945 47805 434979
rect 48053 434945 48087 434979
rect 48237 434945 48271 434979
rect 56793 434945 56827 434979
rect 47869 434809 47903 434843
rect 47961 434809 47995 434843
rect 47593 434741 47627 434775
rect 91477 434265 91511 434299
rect 91661 434265 91695 434299
rect 91845 434265 91879 434299
rect 64061 433381 64095 433415
rect 281365 432157 281399 432191
rect 281632 432089 281666 432123
rect 282745 432021 282779 432055
rect 142261 429505 142295 429539
rect 142445 429505 142479 429539
rect 142353 429369 142387 429403
rect 412281 428417 412315 428451
rect 412373 428417 412407 428451
rect 412005 428349 412039 428383
rect 412557 428281 412591 428315
rect 412097 428213 412131 428247
rect 450553 426717 450587 426751
rect 239137 424541 239171 424575
rect 239321 424541 239355 424575
rect 238953 424473 238987 424507
rect 331413 423521 331447 423555
rect 332057 423521 332091 423555
rect 133705 423453 133739 423487
rect 133888 423453 133922 423487
rect 133981 423453 134015 423487
rect 134119 423453 134153 423487
rect 134257 423453 134291 423487
rect 331137 423453 331171 423487
rect 331320 423453 331354 423487
rect 331505 423453 331539 423487
rect 331689 423453 331723 423487
rect 134349 423317 134383 423351
rect 331781 423317 331815 423351
rect 27537 423113 27571 423147
rect 332057 423113 332091 423147
rect 32045 423045 32079 423079
rect 27445 422977 27479 423011
rect 27997 422977 28031 423011
rect 28273 422977 28307 423011
rect 27629 422909 27663 422943
rect 28365 422909 28399 422943
rect 28365 422773 28399 422807
rect 32045 422773 32079 422807
rect 443929 421277 443963 421311
rect 443662 421209 443696 421243
rect 442549 421141 442583 421175
rect 333989 417537 334023 417571
rect 334081 417537 334115 417571
rect 334357 417469 334391 417503
rect 334265 417401 334299 417435
rect 333805 417333 333839 417367
rect 136557 417129 136591 417163
rect 256525 415497 256559 415531
rect 256893 415429 256927 415463
rect 279709 415429 279743 415463
rect 279249 415361 279283 415395
rect 279341 415361 279375 415395
rect 279893 415361 279927 415395
rect 256985 415293 257019 415327
rect 257077 415293 257111 415327
rect 279065 415293 279099 415327
rect 279617 415293 279651 415327
rect 279525 415225 279559 415259
rect 119629 414749 119663 414783
rect 402693 414273 402727 414307
rect 402437 414205 402471 414239
rect 403817 414069 403851 414103
rect 258917 413865 258951 413899
rect 260297 413661 260331 413695
rect 260030 413593 260064 413627
rect 143825 412777 143859 412811
rect 151461 411893 151495 411927
rect 338405 411485 338439 411519
rect 99665 411009 99699 411043
rect 99849 411009 99883 411043
rect 99941 410873 99975 410907
rect 112545 410601 112579 410635
rect 113005 410601 113039 410635
rect 113097 410465 113131 410499
rect 112729 410397 112763 410431
rect 112821 410397 112855 410431
rect 55321 409921 55355 409955
rect 55505 409921 55539 409955
rect 55689 409921 55723 409955
rect 57805 409513 57839 409547
rect 57161 409377 57195 409411
rect 57253 409377 57287 409411
rect 56885 409309 56919 409343
rect 56977 409309 57011 409343
rect 57805 409241 57839 409275
rect 56701 409173 56735 409207
rect 441813 406045 441847 406079
rect 114109 405569 114143 405603
rect 56609 403189 56643 403223
rect 169953 401693 169987 401727
rect 67189 400673 67223 400707
rect 67097 400605 67131 400639
rect 67373 400605 67407 400639
rect 67465 400605 67499 400639
rect 67649 400469 67683 400503
rect 268945 399925 268979 399959
rect 252937 399517 252971 399551
rect 253121 399381 253155 399415
rect 400045 398429 400079 398463
rect 326537 397749 326571 397783
rect 340797 397477 340831 397511
rect 282653 396253 282687 396287
rect 43085 395777 43119 395811
rect 313749 395573 313783 395607
rect 380541 395233 380575 395267
rect 11805 395165 11839 395199
rect 380725 395165 380759 395199
rect 11989 395029 12023 395063
rect 380909 395029 380943 395063
rect 22845 394825 22879 394859
rect 23397 394825 23431 394859
rect 23029 394689 23063 394723
rect 23397 394689 23431 394723
rect 452117 394145 452151 394179
rect 451933 394077 451967 394111
rect 452025 394009 452059 394043
rect 451565 393941 451599 393975
rect 20545 393397 20579 393431
rect 257077 392309 257111 392343
rect 346777 387617 346811 387651
rect 346869 387617 346903 387651
rect 346501 387549 346535 387583
rect 346593 387549 346627 387583
rect 346317 387413 346351 387447
rect 367753 387073 367787 387107
rect 367845 387073 367879 387107
rect 367477 387005 367511 387039
rect 367569 386937 367603 386971
rect 368029 386869 368063 386903
rect 199393 384761 199427 384795
rect 108313 384693 108347 384727
rect 89453 384489 89487 384523
rect 89269 384353 89303 384387
rect 103345 384285 103379 384319
rect 103437 384285 103471 384319
rect 132601 384285 132635 384319
rect 88809 384217 88843 384251
rect 89085 384149 89119 384183
rect 89177 384149 89211 384183
rect 103529 384149 103563 384183
rect 132417 384149 132451 384183
rect 198013 384149 198047 384183
rect 177037 383945 177071 383979
rect 198013 383877 198047 383911
rect 177221 383809 177255 383843
rect 177313 383809 177347 383843
rect 177589 383809 177623 383843
rect 177497 383673 177531 383707
rect 200589 384149 200623 384183
rect 200037 383877 200071 383911
rect 200589 383877 200623 383911
rect 199945 383809 199979 383843
rect 200405 383809 200439 383843
rect 200129 383741 200163 383775
rect 199393 383605 199427 383639
rect 199577 383605 199611 383639
rect 200405 383605 200439 383639
rect 96353 383197 96387 383231
rect 130393 383197 130427 383231
rect 322305 383197 322339 383231
rect 40785 381021 40819 381055
rect 40518 380953 40552 380987
rect 39405 380885 39439 380919
rect 274465 380409 274499 380443
rect 70685 378845 70719 378879
rect 70869 378845 70903 378879
rect 71881 378845 71915 378879
rect 71329 378777 71363 378811
rect 70593 378709 70627 378743
rect 309701 375785 309735 375819
rect 308321 375649 308355 375683
rect 207581 375581 207615 375615
rect 308566 375513 308600 375547
rect 409429 375105 409463 375139
rect 409521 375037 409555 375071
rect 409613 375037 409647 375071
rect 409061 374901 409095 374935
rect 95617 374697 95651 374731
rect 450461 374697 450495 374731
rect 95985 374561 96019 374595
rect 95801 374493 95835 374527
rect 450645 374493 450679 374527
rect 441997 372317 442031 372351
rect 233709 371841 233743 371875
rect 233801 371637 233835 371671
rect 214757 370141 214791 370175
rect 293693 369053 293727 369087
rect 293785 368917 293819 368951
rect 360577 366537 360611 366571
rect 360393 366401 360427 366435
rect 360209 366333 360243 366367
rect 143457 365449 143491 365483
rect 473737 365449 473771 365483
rect 142997 365381 143031 365415
rect 143181 365381 143215 365415
rect 143365 365313 143399 365347
rect 143457 365313 143491 365347
rect 473645 365313 473679 365347
rect 470425 364701 470459 364735
rect 470670 364633 470704 364667
rect 471805 364565 471839 364599
rect 180441 362593 180475 362627
rect 49893 362525 49927 362559
rect 180257 362525 180291 362559
rect 180073 362457 180107 362491
rect 244381 360349 244415 360383
rect 402805 360349 402839 360383
rect 402989 360349 403023 360383
rect 402897 360213 402931 360247
rect 361497 359873 361531 359907
rect 361681 359669 361715 359703
rect 88349 359329 88383 359363
rect 88165 359261 88199 359295
rect 87981 359125 88015 359159
rect 90649 356745 90683 356779
rect 89525 356609 89559 356643
rect 89269 356541 89303 356575
rect 200037 356065 200071 356099
rect 7481 355997 7515 356031
rect 361589 355997 361623 356031
rect 7389 355861 7423 355895
rect 361405 355861 361439 355895
rect 403725 355317 403759 355351
rect 195069 354365 195103 354399
rect 194425 354229 194459 354263
rect 194149 353821 194183 353855
rect 195897 353821 195931 353855
rect 194793 353753 194827 353787
rect 193689 353685 193723 353719
rect 194609 353413 194643 353447
rect 193597 353345 193631 353379
rect 193689 353345 193723 353379
rect 193965 353345 193999 353379
rect 195437 353345 195471 353379
rect 193413 353277 193447 353311
rect 193873 353277 193907 353311
rect 141065 351645 141099 351679
rect 451473 349469 451507 349503
rect 451565 349333 451599 349367
rect 5365 348585 5399 348619
rect 5365 348449 5399 348483
rect 4721 348381 4755 348415
rect 4905 348381 4939 348415
rect 4997 348381 5031 348415
rect 5090 348381 5124 348415
rect 5273 348381 5307 348415
rect 4629 348245 4663 348279
rect 485421 346817 485455 346851
rect 485605 346817 485639 346851
rect 485513 346613 485547 346647
rect 376217 344437 376251 344471
rect 233341 344233 233375 344267
rect 232697 344097 232731 344131
rect 29561 344029 29595 344063
rect 232881 343893 232915 343927
rect 232973 343893 233007 343927
rect 410993 339677 411027 339711
rect 344753 339201 344787 339235
rect 344569 339133 344603 339167
rect 344937 338997 344971 339031
rect 385141 338113 385175 338147
rect 385233 338113 385267 338147
rect 218989 337705 219023 337739
rect 218805 337569 218839 337603
rect 218713 337501 218747 337535
rect 218989 337433 219023 337467
rect 218529 337365 218563 337399
rect 106114 336005 106148 336039
rect 106381 335937 106415 335971
rect 105001 335733 105035 335767
rect 68201 335325 68235 335359
rect 365821 334645 365855 334679
rect 310897 334305 310931 334339
rect 311725 334305 311759 334339
rect 310621 334237 310655 334271
rect 310805 334237 310839 334271
rect 310990 334234 311024 334268
rect 311173 334237 311207 334271
rect 310529 334101 310563 334135
rect 314485 334169 314519 334203
rect 314669 334237 314703 334271
rect 314761 334237 314795 334271
rect 314669 334033 314703 334067
rect 311725 333965 311759 333999
rect 9597 333149 9631 333183
rect 9873 333149 9907 333183
rect 9321 333081 9355 333115
rect 9505 333013 9539 333047
rect 9689 333013 9723 333047
rect 62221 332605 62255 332639
rect 87797 331381 87831 331415
rect 363521 331177 363555 331211
rect 381553 329545 381587 329579
rect 381645 329545 381679 329579
rect 381461 329409 381495 329443
rect 381829 329409 381863 329443
rect 438317 329409 438351 329443
rect 438501 329409 438535 329443
rect 251189 329341 251223 329375
rect 252385 329341 252419 329375
rect 381277 329273 381311 329307
rect 438409 329205 438443 329239
rect 251189 329001 251223 329035
rect 208501 327709 208535 327743
rect 424057 327369 424091 327403
rect 423965 327233 423999 327267
rect 87061 326621 87095 326655
rect 93317 326145 93351 326179
rect 93501 326145 93535 326179
rect 91569 326009 91603 326043
rect 93685 325941 93719 325975
rect 450553 325533 450587 325567
rect 331597 325057 331631 325091
rect 331781 325057 331815 325091
rect 282285 324989 282319 325023
rect 331873 324853 331907 324887
rect 348433 322677 348467 322711
rect 465457 320161 465491 320195
rect 78965 319413 78999 319447
rect 342269 319073 342303 319107
rect 342002 318937 342036 318971
rect 340889 318869 340923 318903
rect 182097 317373 182131 317407
rect 21281 317237 21315 317271
rect 481833 314313 481867 314347
rect 481741 314177 481775 314211
rect 183385 312137 183419 312171
rect 184498 312069 184532 312103
rect 184765 311933 184799 311967
rect 403357 310709 403391 310743
rect 426817 308737 426851 308771
rect 426909 308737 426943 308771
rect 426449 308669 426483 308703
rect 426541 308669 426575 308703
rect 427093 308601 427127 308635
rect 426449 308533 426483 308567
rect 426633 308533 426667 308567
rect 140697 307105 140731 307139
rect 140789 306969 140823 307003
rect 140881 306901 140915 306935
rect 141249 306901 141283 306935
rect 187433 306357 187467 306391
rect 22109 306153 22143 306187
rect 21465 306017 21499 306051
rect 21649 306017 21683 306051
rect 21741 305813 21775 305847
rect 49893 304861 49927 304895
rect 50077 304861 50111 304895
rect 5834 304453 5868 304487
rect 50322 304793 50356 304827
rect 51457 304725 51491 304759
rect 6101 304317 6135 304351
rect 49893 304317 49927 304351
rect 4721 304181 4755 304215
rect 325801 303093 325835 303127
rect 262505 301597 262539 301631
rect 262238 301529 262272 301563
rect 261125 301461 261159 301495
rect 341073 301121 341107 301155
rect 340889 301053 340923 301087
rect 341257 300917 341291 300951
rect 46489 298333 46523 298367
rect 414213 296157 414247 296191
rect 414397 296157 414431 296191
rect 414581 296021 414615 296055
rect 112821 295817 112855 295851
rect 111993 295681 112027 295715
rect 112176 295681 112210 295715
rect 112545 295681 112579 295715
rect 112269 295613 112303 295647
rect 112361 295613 112395 295647
rect 112821 295613 112855 295647
rect 112637 295477 112671 295511
rect 104541 293981 104575 294015
rect 274741 293301 274775 293335
rect 84209 292893 84243 292927
rect 138193 292417 138227 292451
rect 137937 292349 137971 292383
rect 139317 292213 139351 292247
rect 340889 291329 340923 291363
rect 341258 291329 341292 291363
rect 341441 291329 341475 291363
rect 341073 291261 341107 291295
rect 341165 291261 341199 291295
rect 340705 291193 340739 291227
rect 92949 288065 92983 288099
rect 93133 288065 93167 288099
rect 92765 287861 92799 287895
rect 273637 286977 273671 287011
rect 273821 286977 273855 287011
rect 274005 286841 274039 286875
rect 244473 283849 244507 283883
rect 243349 283713 243383 283747
rect 297557 283713 297591 283747
rect 243093 283645 243127 283679
rect 297281 283645 297315 283679
rect 296085 283305 296119 283339
rect 483029 283305 483063 283339
rect 297649 283169 297683 283203
rect 296269 283101 296303 283135
rect 296729 283101 296763 283135
rect 296269 282761 296303 282795
rect 296085 282625 296119 282659
rect 296913 282625 296947 282659
rect 297925 282557 297959 282591
rect 16865 282013 16899 282047
rect 84577 281333 84611 281367
rect 329757 280449 329791 280483
rect 329665 280245 329699 280279
rect 264612 279429 264646 279463
rect 264345 279361 264379 279395
rect 265725 279157 265759 279191
rect 176945 277865 176979 277899
rect 248705 276097 248739 276131
rect 248613 276029 248647 276063
rect 158729 273921 158763 273955
rect 158912 273921 158946 273955
rect 159097 273921 159131 273955
rect 159281 273921 159315 273955
rect 159005 273853 159039 273887
rect 159373 273717 159407 273751
rect 229109 273309 229143 273343
rect 420561 272629 420595 272663
rect 373273 271269 373307 271303
rect 373089 271133 373123 271167
rect 373733 271133 373767 271167
rect 374929 271065 374963 271099
rect 375297 271065 375331 271099
rect 373825 270793 373859 270827
rect 374285 270657 374319 270691
rect 375297 270657 375331 270691
rect 92305 270249 92339 270283
rect 92489 270045 92523 270079
rect 228741 267869 228775 267903
rect 228925 267869 228959 267903
rect 229109 267733 229143 267767
rect 367293 266781 367327 266815
rect 367477 266781 367511 266815
rect 486985 266781 487019 266815
rect 486718 266713 486752 266747
rect 367109 266645 367143 266679
rect 485605 266645 485639 266679
rect 36369 266305 36403 266339
rect 353401 265761 353435 265795
rect 442273 265693 442307 265727
rect 78128 264129 78162 264163
rect 77861 264061 77895 264095
rect 79241 263925 79275 263959
rect 98745 263925 98779 263959
rect 207397 262565 207431 262599
rect 207121 262429 207155 262463
rect 207397 262429 207431 262463
rect 125893 261001 125927 261035
rect 126069 261001 126103 261035
rect 125517 260933 125551 260967
rect 125333 260865 125367 260899
rect 125609 260865 125643 260899
rect 125753 260865 125787 260899
rect 126069 260865 126103 260899
rect 317797 260253 317831 260287
rect 317705 260117 317739 260151
rect 180717 259233 180751 259267
rect 60013 259165 60047 259199
rect 180901 259097 180935 259131
rect 180809 259029 180843 259063
rect 181269 259029 181303 259063
rect 483765 257601 483799 257635
rect 483581 257533 483615 257567
rect 483949 257397 483983 257431
rect 470517 256989 470551 257023
rect 470609 256853 470643 256887
rect 299397 256649 299431 256683
rect 299121 256513 299155 256547
rect 299213 256513 299247 256547
rect 298845 256445 298879 256479
rect 298937 256309 298971 256343
rect 220553 254881 220587 254915
rect 396641 254813 396675 254847
rect 220286 254745 220320 254779
rect 219173 254677 219207 254711
rect 380633 254133 380667 254167
rect 117605 252841 117639 252875
rect 139041 252773 139075 252807
rect 117789 252637 117823 252671
rect 117973 252637 118007 252671
rect 444021 252161 444055 252195
rect 444113 252093 444147 252127
rect 444205 252093 444239 252127
rect 443653 251957 443687 251991
rect 231205 251073 231239 251107
rect 230949 251005 230983 251039
rect 232329 250937 232363 250971
rect 303169 249985 303203 250019
rect 302985 249781 303019 249815
rect 315129 248693 315163 248727
rect 115213 244341 115247 244375
rect 315773 240873 315807 240907
rect 468033 240873 468067 240907
rect 467389 240601 467423 240635
rect 467849 240601 467883 240635
rect 467665 240533 467699 240567
rect 467757 240533 467791 240567
rect 20545 237541 20579 237575
rect 430957 237541 430991 237575
rect 20361 237405 20395 237439
rect 430773 237405 430807 237439
rect 61117 236317 61151 236351
rect 342545 236317 342579 236351
rect 61384 236249 61418 236283
rect 342278 236249 342312 236283
rect 62497 236181 62531 236215
rect 341165 236181 341199 236215
rect 240333 232441 240367 232475
rect 216229 231489 216263 231523
rect 418537 231013 418571 231047
rect 419089 230945 419123 230979
rect 418905 230809 418939 230843
rect 418997 230741 419031 230775
rect 153393 229789 153427 229823
rect 153485 229789 153519 229823
rect 167837 228361 167871 228395
rect 167469 228225 167503 228259
rect 167193 228157 167227 228191
rect 167377 228157 167411 228191
rect 292221 228021 292255 228055
rect 137201 227681 137235 227715
rect 136465 227613 136499 227647
rect 136741 227273 136775 227307
rect 135637 227137 135671 227171
rect 135913 227137 135947 227171
rect 136006 227137 136040 227171
rect 136189 227137 136223 227171
rect 135821 227069 135855 227103
rect 137201 227069 137235 227103
rect 135545 226933 135579 226967
rect 347053 225641 347087 225675
rect 290289 224961 290323 224995
rect 289829 224757 289863 224791
rect 100861 224553 100895 224587
rect 290013 224553 290047 224587
rect 289461 224417 289495 224451
rect 100953 224349 100987 224383
rect 289553 224213 289587 224247
rect 289645 224213 289679 224247
rect 265725 223533 265759 223567
rect 227913 223465 227947 223499
rect 265725 223329 265759 223363
rect 260481 223261 260515 223295
rect 260849 223261 260883 223295
rect 260665 223125 260699 223159
rect 260849 223125 260883 223159
rect 79793 220745 79827 220779
rect 97089 220745 97123 220779
rect 123401 220745 123435 220779
rect 131865 220745 131899 220779
rect 164157 220745 164191 220779
rect 205649 220745 205683 220779
rect 128461 220677 128495 220711
rect 129657 220677 129691 220711
rect 259285 220677 259319 220711
rect 266645 220677 266679 220711
rect 50077 220609 50111 220643
rect 75745 220609 75779 220643
rect 75837 220609 75871 220643
rect 79425 220609 79459 220643
rect 96721 220609 96755 220643
rect 123493 220609 123527 220643
rect 124137 220609 124171 220643
rect 55045 220473 55079 220507
rect 75653 220473 75687 220507
rect 78965 220541 78999 220575
rect 79149 220541 79183 220575
rect 79333 220541 79367 220575
rect 96169 220541 96203 220575
rect 96445 220541 96479 220575
rect 96629 220541 96663 220575
rect 97181 220541 97215 220575
rect 49985 220405 50019 220439
rect 75837 220405 75871 220439
rect 77769 220405 77803 220439
rect 78965 220405 78999 220439
rect 96169 220405 96203 220439
rect 97181 220405 97215 220439
rect 124137 219861 124171 219895
rect 128369 220609 128403 220643
rect 11805 219521 11839 219555
rect 9505 219045 9539 219079
rect 12817 219521 12851 219555
rect 16221 219521 16255 219555
rect 17233 219521 17267 219555
rect 96077 219521 96111 219555
rect 53757 219453 53791 219487
rect 22937 219317 22971 219351
rect 22937 218773 22971 218807
rect 78137 219317 78171 219351
rect 78137 218841 78171 218875
rect 96077 218841 96111 218875
rect 114385 219317 114419 219351
rect 53757 218773 53791 218807
rect 17233 218637 17267 218671
rect 16221 218569 16255 218603
rect 12817 218501 12851 218535
rect 11805 218433 11839 218467
rect 128369 218977 128403 219011
rect 129565 220609 129599 220643
rect 132989 220609 133023 220643
rect 133797 220609 133831 220643
rect 163044 220609 163078 220643
rect 167101 220609 167135 220643
rect 178325 220609 178359 220643
rect 205005 220609 205039 220643
rect 205188 220609 205222 220643
rect 205281 220609 205315 220643
rect 205557 220609 205591 220643
rect 235273 220609 235307 220643
rect 257445 220609 257479 220643
rect 257537 220609 257571 220643
rect 257997 220609 258031 220643
rect 259096 220609 259130 220643
rect 259193 220609 259227 220643
rect 259468 220609 259502 220643
rect 259561 220609 259595 220643
rect 266205 220609 266239 220643
rect 129105 220541 129139 220575
rect 129381 220541 129415 220575
rect 133245 220541 133279 220575
rect 130025 220405 130059 220439
rect 162777 220541 162811 220575
rect 133797 220133 133831 220167
rect 205373 220541 205407 220575
rect 257169 220541 257203 220575
rect 257261 220541 257295 220575
rect 204821 220473 204855 220507
rect 178049 220405 178083 220439
rect 178417 220405 178451 220439
rect 178049 220065 178083 220099
rect 167101 219997 167135 220031
rect 129105 219929 129139 219963
rect 257721 220405 257755 220439
rect 266461 220541 266495 220575
rect 258089 220405 258123 220439
rect 258917 220405 258951 220439
rect 265081 220405 265115 220439
rect 258089 220065 258123 220099
rect 257997 219929 258031 219963
rect 204821 219861 204855 219895
rect 267013 220609 267047 220643
rect 287621 220609 287655 220643
rect 288265 220609 288299 220643
rect 267013 220065 267047 220099
rect 272441 220541 272475 220575
rect 272533 220541 272567 220575
rect 272533 220337 272567 220371
rect 272441 220065 272475 220099
rect 266645 219861 266679 219895
rect 266737 219861 266771 219895
rect 254961 219793 254995 219827
rect 254961 219657 254995 219691
rect 266737 219657 266771 219691
rect 287621 219453 287655 219487
rect 128461 218909 128495 218943
rect 232973 219317 233007 219351
rect 232973 218705 233007 218739
rect 248337 219317 248371 219351
rect 248337 218705 248371 218739
rect 114385 218229 114419 218263
rect 345857 218229 345891 218263
rect 9505 217685 9539 217719
rect 370973 216937 371007 216971
rect 370881 216869 370915 216903
rect 370973 216801 371007 216835
rect 371249 216801 371283 216835
rect 370881 216733 370915 216767
rect 371157 216733 371191 216767
rect 371433 216733 371467 216767
rect 371525 216733 371559 216767
rect 371709 216665 371743 216699
rect 310069 210409 310103 210443
rect 3249 209525 3283 209559
rect 9505 203881 9539 203915
rect 9321 203677 9355 203711
rect 310069 202113 310103 202147
rect 310345 201909 310379 201943
rect 310529 201909 310563 201943
rect 413753 200821 413787 200855
rect 483857 199937 483891 199971
rect 450553 195381 450587 195415
rect 397469 194973 397503 195007
rect 310344 183617 310378 183651
rect 310437 183617 310471 183651
rect 310529 183617 310563 183651
rect 310713 183617 310747 183651
rect 310069 183549 310103 183583
rect 406393 179741 406427 179775
rect 407589 179741 407623 179775
rect 406853 179605 406887 179639
rect 407405 179605 407439 179639
rect 310161 178313 310195 178347
rect 310345 178177 310379 178211
rect 310437 178177 310471 178211
rect 310713 178109 310747 178143
rect 310621 178041 310655 178075
rect 310253 176137 310287 176171
rect 336197 176137 336231 176171
rect 336565 176137 336599 176171
rect 336105 176069 336139 176103
rect 310069 176001 310103 176035
rect 335921 175933 335955 175967
rect 337025 175933 337059 175967
rect 337485 175797 337519 175831
rect 3617 170153 3651 170187
rect 4997 170017 5031 170051
rect 4741 169949 4775 169983
rect 380725 161993 380759 162027
rect 381093 161993 381127 162027
rect 385417 161925 385451 161959
rect 385049 161857 385083 161891
rect 385233 161857 385267 161891
rect 385601 161857 385635 161891
rect 385785 161857 385819 161891
rect 381185 161789 381219 161823
rect 381369 161789 381403 161823
rect 414857 161653 414891 161687
rect 466009 161653 466043 161687
rect 8125 157097 8159 157131
rect 484225 157097 484259 157131
rect 8217 156893 8251 156927
rect 321477 152609 321511 152643
rect 323593 152609 323627 152643
rect 322029 152405 322063 152439
rect 322489 152405 322523 152439
rect 323041 152405 323075 152439
rect 322305 152133 322339 152167
rect 321661 152065 321695 152099
rect 321753 152065 321787 152099
rect 322029 152065 322063 152099
rect 427277 152065 427311 152099
rect 321937 151997 321971 152031
rect 321477 151861 321511 151895
rect 357357 148189 357391 148223
rect 315497 147509 315531 147543
rect 9505 145333 9539 145367
rect 9597 145129 9631 145163
rect 389373 143157 389407 143191
rect 454969 142749 455003 142783
rect 9597 142137 9631 142171
rect 9781 142273 9815 142307
rect 9413 136425 9447 136459
rect 457729 142137 457763 142171
rect 416145 140573 416179 140607
rect 416412 140505 416446 140539
rect 417525 140437 417559 140471
rect 7481 136357 7515 136391
rect 9781 136357 9815 136391
rect 9321 136221 9355 136255
rect 7297 135337 7331 135371
rect 7481 135337 7515 135371
rect 8769 133093 8803 133127
rect 9229 133025 9263 133059
rect 8953 132957 8987 132991
rect 9137 132957 9171 132991
rect 9322 132957 9356 132991
rect 9505 132957 9539 132991
rect 355977 132957 356011 132991
rect 356713 128605 356747 128639
rect 4537 127517 4571 127551
rect 4721 127381 4755 127415
rect 383669 126429 383703 126463
rect 477785 126089 477819 126123
rect 477693 125953 477727 125987
rect 428933 124865 428967 124899
rect 429209 124865 429243 124899
rect 429301 124865 429335 124899
rect 429485 124729 429519 124763
rect 429025 124661 429059 124695
rect 310253 123573 310287 123607
rect 366833 123369 366867 123403
rect 366741 123233 366775 123267
rect 367017 123165 367051 123199
rect 367109 123165 367143 123199
rect 367293 123029 367327 123063
rect 299673 120853 299707 120887
rect 248889 120785 248923 120819
rect 248889 120649 248923 120683
rect 299673 120649 299707 120683
rect 239597 120037 239631 120071
rect 156613 119901 156647 119935
rect 80989 119833 81023 119867
rect 75745 119765 75779 119799
rect 34989 119425 35023 119459
rect 35173 119425 35207 119459
rect 35358 119425 35392 119459
rect 35541 119425 35575 119459
rect 35725 119425 35759 119459
rect 38761 119425 38795 119459
rect 61209 119425 61243 119459
rect 63693 119425 63727 119459
rect 63877 119425 63911 119459
rect 64061 119425 64095 119459
rect 35265 119357 35299 119391
rect 33517 119221 33551 119255
rect 34897 119221 34931 119255
rect 75561 119289 75595 119323
rect 75745 119289 75779 119323
rect 145297 119425 145331 119459
rect 145481 119425 145515 119459
rect 145665 119425 145699 119459
rect 80989 119289 81023 119323
rect 81357 119289 81391 119323
rect 38853 119221 38887 119255
rect 102701 119221 102735 119255
rect 34621 119017 34655 119051
rect 35725 119017 35759 119051
rect 43821 118949 43855 118983
rect 35081 118881 35115 118915
rect 34805 118813 34839 118847
rect 34897 118813 34931 118847
rect 35173 118813 35207 118847
rect 166273 119901 166307 119935
rect 162164 119493 162198 119527
rect 233893 119901 233927 119935
rect 239229 119901 239263 119935
rect 239321 119901 239355 119935
rect 233893 119629 233927 119663
rect 215585 119425 215619 119459
rect 215769 119425 215803 119459
rect 215861 119425 215895 119459
rect 216137 119425 216171 119459
rect 233893 119425 233927 119459
rect 238769 119425 238803 119459
rect 238861 119425 238895 119459
rect 156613 119357 156647 119391
rect 162409 119357 162443 119391
rect 166273 119357 166307 119391
rect 214481 119357 214515 119391
rect 216045 119357 216079 119391
rect 233341 119357 233375 119391
rect 234077 119357 234111 119391
rect 239137 119357 239171 119391
rect 239229 119357 239263 119391
rect 239505 119357 239539 119391
rect 145757 119289 145791 119323
rect 161029 119221 161063 119255
rect 172713 119221 172747 119255
rect 214481 118949 214515 118983
rect 216321 119289 216355 119323
rect 233341 119221 233375 119255
rect 238309 119289 238343 119323
rect 216321 118949 216355 118983
rect 238585 119221 238619 119255
rect 239045 119221 239079 119255
rect 289829 119969 289863 120003
rect 258641 119697 258675 119731
rect 248521 119629 248555 119663
rect 248429 119357 248463 119391
rect 253121 119493 253155 119527
rect 254225 119425 254259 119459
rect 254317 119425 254351 119459
rect 255237 119425 255271 119459
rect 253121 119289 253155 119323
rect 248337 119221 248371 119255
rect 239321 119153 239355 119187
rect 239597 119153 239631 119187
rect 253949 119153 253983 119187
rect 239321 118813 239355 118847
rect 248521 119017 248555 119051
rect 248521 118813 248555 118847
rect 254501 119085 254535 119119
rect 254225 118813 254259 118847
rect 258641 119289 258675 119323
rect 258733 119425 258767 119459
rect 289921 119969 289955 120003
rect 291853 119969 291887 120003
rect 290013 119697 290047 119731
rect 290749 119697 290783 119731
rect 289921 119629 289955 119663
rect 291853 119629 291887 119663
rect 291945 119969 291979 120003
rect 307677 119765 307711 119799
rect 308229 119697 308263 119731
rect 291945 119493 291979 119527
rect 290289 119425 290323 119459
rect 290565 119425 290599 119459
rect 289829 119357 289863 119391
rect 290197 119357 290231 119391
rect 258733 119221 258767 119255
rect 301605 119289 301639 119323
rect 255237 118881 255271 118915
rect 258917 119085 258951 119119
rect 238309 118745 238343 118779
rect 253949 118745 253983 118779
rect 291945 119085 291979 119119
rect 291853 118881 291887 118915
rect 289277 118813 289311 118847
rect 289461 118813 289495 118847
rect 258917 118745 258951 118779
rect 291853 118745 291887 118779
rect 297925 119085 297959 119119
rect 301605 119085 301639 119119
rect 307677 119289 307711 119323
rect 308045 119289 308079 119323
rect 297925 118881 297959 118915
rect 308229 119085 308263 119119
rect 307677 118813 307711 118847
rect 291945 118745 291979 118779
rect 307493 118745 307527 118779
rect 145297 118677 145331 118711
rect 451390 117249 451424 117283
rect 451657 117249 451691 117283
rect 450277 117045 450311 117079
rect 485237 117045 485271 117079
rect 224325 116637 224359 116671
rect 209513 115753 209547 115787
rect 209881 115617 209915 115651
rect 209697 115549 209731 115583
rect 440341 114869 440375 114903
rect 32597 113985 32631 114019
rect 32505 113849 32539 113883
rect 69213 113373 69247 113407
rect 69397 113373 69431 113407
rect 69029 113237 69063 113271
rect 328561 112217 328595 112251
rect 328285 112149 328319 112183
rect 327733 111945 327767 111979
rect 327273 111809 327307 111843
rect 327365 111809 327399 111843
rect 328561 111809 328595 111843
rect 329573 111809 329607 111843
rect 329757 111809 329791 111843
rect 132049 111741 132083 111775
rect 84025 111401 84059 111435
rect 28641 111129 28675 111163
rect 82829 110857 82863 110891
rect 83105 110857 83139 110891
rect 83473 110857 83507 110891
rect 28457 110721 28491 110755
rect 28641 110721 28675 110755
rect 50537 110721 50571 110755
rect 50997 110721 51031 110755
rect 18981 110653 19015 110687
rect 83565 110721 83599 110755
rect 106289 111061 106323 111095
rect 96905 110721 96939 110755
rect 82829 110653 82863 110687
rect 83749 110653 83783 110687
rect 84025 110653 84059 110687
rect 108313 111061 108347 111095
rect 106473 110721 106507 110755
rect 106740 110721 106774 110755
rect 106289 110653 106323 110687
rect 108313 110653 108347 110687
rect 108405 111061 108439 111095
rect 50997 110585 51031 110619
rect 326813 111741 326847 111775
rect 327181 111741 327215 111775
rect 327917 111741 327951 111775
rect 179061 111673 179095 111707
rect 166273 111469 166307 111503
rect 170505 111469 170539 111503
rect 173817 111469 173851 111503
rect 178969 111469 179003 111503
rect 173817 111333 173851 111367
rect 173909 111333 173943 111367
rect 183385 111673 183419 111707
rect 179061 111333 179095 111367
rect 179153 111333 179187 111367
rect 178969 111197 179003 111231
rect 179521 111197 179555 111231
rect 179613 111197 179647 111231
rect 182005 111197 182039 111231
rect 182925 111197 182959 111231
rect 183109 111197 183143 111231
rect 179153 111129 179187 111163
rect 179981 111129 180015 111163
rect 173909 111061 173943 111095
rect 179337 111061 179371 111095
rect 178693 110789 178727 110823
rect 166273 110721 166307 110755
rect 168113 110721 168147 110755
rect 168297 110721 168331 110755
rect 170321 110721 170355 110755
rect 170413 110721 170447 110755
rect 170505 110721 170539 110755
rect 178601 110721 178635 110755
rect 168113 110585 168147 110619
rect 101045 110517 101079 110551
rect 107853 110517 107887 110551
rect 108405 110517 108439 110551
rect 131497 110517 131531 110551
rect 132049 110517 132083 110551
rect 137201 110517 137235 110551
rect 170229 110517 170263 110551
rect 170413 110517 170447 110551
rect 181085 110789 181119 110823
rect 180634 110721 180668 110755
rect 180901 110653 180935 110687
rect 179521 110517 179555 110551
rect 178693 110245 178727 110279
rect 221657 111537 221691 111571
rect 183293 111061 183327 111095
rect 183385 111061 183419 111095
rect 187801 111469 187835 111503
rect 182649 110721 182683 110755
rect 182741 110721 182775 110755
rect 183109 110721 183143 110755
rect 183201 110721 183235 110755
rect 181545 110653 181579 110687
rect 182097 110653 182131 110687
rect 181085 110245 181119 110279
rect 178601 110177 178635 110211
rect 194885 111469 194919 111503
rect 191021 111333 191055 111367
rect 187801 110925 187835 110959
rect 190101 111197 190135 111231
rect 190929 111197 190963 111231
rect 191021 111197 191055 111231
rect 190101 110857 190135 110891
rect 183293 110653 183327 110687
rect 194885 110857 194919 110891
rect 202521 111333 202555 111367
rect 194425 110721 194459 110755
rect 194563 110721 194597 110755
rect 191021 110585 191055 110619
rect 194609 110585 194643 110619
rect 190469 110517 190503 110551
rect 212641 111197 212675 111231
rect 212641 110789 212675 110823
rect 222761 111401 222795 111435
rect 214481 110721 214515 110755
rect 214665 110721 214699 110755
rect 221749 110721 221783 110755
rect 221838 110721 221872 110755
rect 222024 110721 222058 110755
rect 222209 110721 222243 110755
rect 222393 110721 222427 110755
rect 221657 110653 221691 110687
rect 222112 110653 222146 110687
rect 202705 110517 202739 110551
rect 214389 110517 214423 110551
rect 202521 110449 202555 110483
rect 222945 111197 222979 111231
rect 273637 111197 273671 111231
rect 326813 111197 326847 111231
rect 272441 111129 272475 111163
rect 272441 110925 272475 110959
rect 274097 111129 274131 111163
rect 274097 110925 274131 110959
rect 274189 111129 274223 111163
rect 273545 110857 273579 110891
rect 222945 110789 222979 110823
rect 328009 111741 328043 111775
rect 480637 111605 480671 111639
rect 328009 111197 328043 111231
rect 328745 111197 328779 111231
rect 329757 111197 329791 111231
rect 327917 111061 327951 111095
rect 328285 111061 328319 111095
rect 222761 110585 222795 110619
rect 224969 110653 225003 110687
rect 222485 110517 222519 110551
rect 224969 110449 225003 110483
rect 225245 110653 225279 110687
rect 273637 110653 273671 110687
rect 273821 110653 273855 110687
rect 274189 110653 274223 110687
rect 282101 110925 282135 110959
rect 282101 110653 282135 110687
rect 286425 110925 286459 110959
rect 286425 110653 286459 110687
rect 286517 110653 286551 110687
rect 221657 110245 221691 110279
rect 273177 110517 273211 110551
rect 286241 110517 286275 110551
rect 286517 110449 286551 110483
rect 225245 110245 225279 110279
rect 183201 110177 183235 110211
rect 453037 109157 453071 109191
rect 453221 109021 453255 109055
rect 419365 107933 419399 107967
rect 419549 107933 419583 107967
rect 496369 107933 496403 107967
rect 419733 107797 419767 107831
rect 456993 106301 457027 106335
rect 368397 105417 368431 105451
rect 368581 105281 368615 105315
rect 3525 101065 3559 101099
rect 3709 101065 3743 101099
rect 3617 100997 3651 101031
rect 3893 100793 3927 100827
rect 3341 100725 3375 100759
rect 487905 100725 487939 100759
rect 458189 99229 458223 99263
rect 457922 99161 457956 99195
rect 456809 99093 456843 99127
rect 438838 90117 438872 90151
rect 438593 90049 438627 90083
rect 439973 89845 440007 89879
rect 380909 85765 380943 85799
rect 382105 85697 382139 85731
rect 380909 85629 380943 85663
rect 382197 85629 382231 85663
rect 382289 85629 382323 85663
rect 381737 85561 381771 85595
rect 310161 84745 310195 84779
rect 310253 84609 310287 84643
rect 8861 79849 8895 79883
rect 9229 79713 9263 79747
rect 8953 79645 8987 79679
rect 9137 79645 9171 79679
rect 9322 79645 9356 79679
rect 9505 79645 9539 79679
rect 443101 79237 443135 79271
rect 442917 79169 442951 79203
rect 443193 78965 443227 78999
rect 337761 78625 337795 78659
rect 338221 78625 338255 78659
rect 469873 78625 469907 78659
rect 337669 78557 337703 78591
rect 337945 78557 337979 78591
rect 338037 78557 338071 78591
rect 339279 78557 339313 78591
rect 469597 78557 469631 78591
rect 469689 78557 469723 78591
rect 469965 78557 469999 78591
rect 338865 78421 338899 78455
rect 469413 78421 469447 78455
rect 429853 75497 429887 75531
rect 429669 75293 429703 75327
rect 378793 72641 378827 72675
rect 378885 72573 378919 72607
rect 378977 72573 379011 72607
rect 378425 72437 378459 72471
rect 496461 72233 496495 72267
rect 394157 70397 394191 70431
rect 310069 67337 310103 67371
rect 310253 67201 310287 67235
rect 360301 66589 360335 66623
rect 360117 66453 360151 66487
rect 9321 66113 9355 66147
rect 9505 65977 9539 66011
rect 493885 65501 493919 65535
rect 477325 63733 477359 63767
rect 445953 61217 445987 61251
rect 446045 61217 446079 61251
rect 445677 61149 445711 61183
rect 445769 61149 445803 61183
rect 445493 61013 445527 61047
rect 372537 59585 372571 59619
rect 372721 59585 372755 59619
rect 406117 59585 406151 59619
rect 406301 59585 406335 59619
rect 406393 59585 406427 59619
rect 406486 59585 406520 59619
rect 406761 59449 406795 59483
rect 372353 59381 372387 59415
rect 7849 58497 7883 58531
rect 421941 57409 421975 57443
rect 422033 57205 422067 57239
rect 9505 54825 9539 54859
rect 401241 54621 401275 54655
rect 401149 54485 401183 54519
rect 310069 50269 310103 50303
rect 310161 50133 310195 50167
rect 310069 48229 310103 48263
rect 463893 48093 463927 48127
rect 346133 46325 346167 46359
rect 340613 46053 340647 46087
rect 340153 45985 340187 46019
rect 340245 45985 340279 46019
rect 339969 45917 340003 45951
rect 340338 45917 340372 45951
rect 340521 45917 340555 45951
rect 340613 45917 340647 45951
rect 498209 45917 498243 45951
rect 339877 45781 339911 45815
rect 310069 45033 310103 45067
rect 310621 44897 310655 44931
rect 310437 44829 310471 44863
rect 310529 44693 310563 44727
rect 310253 43061 310287 43095
rect 8300 42245 8334 42279
rect 8033 42109 8067 42143
rect 9413 41973 9447 42007
rect 366833 39797 366867 39831
rect 418261 37825 418295 37859
rect 418353 37757 418387 37791
rect 418445 37757 418479 37791
rect 310253 37621 310287 37655
rect 417893 37621 417927 37655
rect 342545 36329 342579 36363
rect 343925 36125 343959 36159
rect 343680 36057 343714 36091
rect 390937 35241 390971 35275
rect 392050 35037 392084 35071
rect 392317 35037 392351 35071
rect 392501 35037 392535 35071
rect 371801 34697 371835 34731
rect 372914 34561 372948 34595
rect 373181 34561 373215 34595
rect 392501 34493 392535 34527
rect 399493 31977 399527 32011
rect 417525 31433 417559 31467
rect 416614 31365 416648 31399
rect 418638 31297 418672 31331
rect 418905 31297 418939 31331
rect 416881 31229 416915 31263
rect 415501 31093 415535 31127
rect 408509 30685 408543 30719
rect 320465 30277 320499 30311
rect 320373 30209 320407 30243
rect 376033 27421 376067 27455
rect 9321 25857 9355 25891
rect 9505 25789 9539 25823
rect 9137 25653 9171 25687
rect 310161 25313 310195 25347
rect 310345 25313 310379 25347
rect 310437 25245 310471 25279
rect 310805 25109 310839 25143
rect 456073 16065 456107 16099
rect 455889 15861 455923 15895
rect 335427 15453 335461 15487
rect 335552 15431 335586 15465
rect 335645 15453 335679 15487
rect 335829 15453 335863 15487
rect 496369 15453 496403 15487
rect 335185 15385 335219 15419
rect 496461 15317 496495 15351
rect 479257 14025 479291 14059
rect 479349 13957 479383 13991
rect 478797 13821 478831 13855
rect 479441 13821 479475 13855
rect 478797 13685 478831 13719
rect 478889 13685 478923 13719
rect 344661 12393 344695 12427
rect 278145 9877 278179 9911
rect 78229 9673 78263 9707
rect 151277 9673 151311 9707
rect 185409 9673 185443 9707
rect 35357 9537 35391 9571
rect 35725 9537 35759 9571
rect 65349 9537 65383 9571
rect 66177 9537 66211 9571
rect 77125 9537 77159 9571
rect 77217 9537 77251 9571
rect 77493 9537 77527 9571
rect 77861 9537 77895 9571
rect 78045 9537 78079 9571
rect 78413 9537 78447 9571
rect 78873 9537 78907 9571
rect 79057 9537 79091 9571
rect 88441 9537 88475 9571
rect 88625 9537 88659 9571
rect 95157 9537 95191 9571
rect 115857 9537 115891 9571
rect 116501 9537 116535 9571
rect 116593 9537 116627 9571
rect 116777 9537 116811 9571
rect 147965 9537 147999 9571
rect 148057 9537 148091 9571
rect 151001 9537 151035 9571
rect 151093 9537 151127 9571
rect 151737 9537 151771 9571
rect 152565 9537 152599 9571
rect 152749 9537 152783 9571
rect 152933 9537 152967 9571
rect 168932 9537 168966 9571
rect 35541 9333 35575 9367
rect 65165 9401 65199 9435
rect 35725 9129 35759 9163
rect 76757 9401 76791 9435
rect 77033 9401 77067 9435
rect 72249 9333 72283 9367
rect 79241 9469 79275 9503
rect 88349 9401 88383 9435
rect 116041 9469 116075 9503
rect 116225 9469 116259 9503
rect 121469 9469 121503 9503
rect 138029 9469 138063 9503
rect 138397 9469 138431 9503
rect 148333 9469 148367 9503
rect 148977 9469 149011 9503
rect 77953 9333 77987 9367
rect 98837 9333 98871 9367
rect 111717 9333 111751 9367
rect 115857 9333 115891 9367
rect 115949 9333 115983 9367
rect 115949 8925 115983 8959
rect 116317 9333 116351 9367
rect 120089 9333 120123 9367
rect 121193 9333 121227 9367
rect 121469 9333 121503 9367
rect 116041 8789 116075 8823
rect 142169 9401 142203 9435
rect 147781 9333 147815 9367
rect 148241 9333 148275 9367
rect 148517 9333 148551 9367
rect 142169 9265 142203 9299
rect 138397 8993 138431 9027
rect 120089 8721 120123 8755
rect 77493 8585 77527 8619
rect 76757 8517 76791 8551
rect 150541 9469 150575 9503
rect 150725 9469 150759 9503
rect 150449 9333 150483 9367
rect 150357 9061 150391 9095
rect 150357 8857 150391 8891
rect 148977 8721 149011 8755
rect 152473 9401 152507 9435
rect 150817 9333 150851 9367
rect 151737 9333 151771 9367
rect 150541 9061 150575 9095
rect 150449 8653 150483 8687
rect 153025 9469 153059 9503
rect 168665 9469 168699 9503
rect 161489 9333 161523 9367
rect 154037 9197 154071 9231
rect 161489 9197 161523 9231
rect 168389 9333 168423 9367
rect 170045 9333 170079 9367
rect 170321 9333 170355 9367
rect 154037 9061 154071 9095
rect 153025 8857 153059 8891
rect 153117 8857 153151 8891
rect 152933 8653 152967 8687
rect 148517 8381 148551 8415
rect 168481 9197 168515 9231
rect 168481 9061 168515 9095
rect 186237 9673 186271 9707
rect 239965 9673 239999 9707
rect 248153 9673 248187 9707
rect 270969 9673 271003 9707
rect 271521 9673 271555 9707
rect 277777 9673 277811 9707
rect 278053 9673 278087 9707
rect 185501 9537 185535 9571
rect 185501 9333 185535 9367
rect 185777 9333 185811 9367
rect 185409 9265 185443 9299
rect 191205 9537 191239 9571
rect 239873 9537 239907 9571
rect 240057 9537 240091 9571
rect 241529 9537 241563 9571
rect 244565 9537 244599 9571
rect 244657 9537 244691 9571
rect 244841 9537 244875 9571
rect 245577 9537 245611 9571
rect 191205 9333 191239 9367
rect 233893 9401 233927 9435
rect 186237 9265 186271 9299
rect 170321 9061 170355 9095
rect 153117 8381 153151 8415
rect 168297 8585 168331 8619
rect 168389 8585 168423 8619
rect 168297 8381 168331 8415
rect 171793 9197 171827 9231
rect 233893 9197 233927 9231
rect 233801 9061 233835 9095
rect 244289 9469 244323 9503
rect 244381 9469 244415 9503
rect 241529 8857 241563 8891
rect 243461 9401 243495 9435
rect 243461 8857 243495 8891
rect 245117 9401 245151 9435
rect 171793 8585 171827 8619
rect 230397 8789 230431 8823
rect 233801 8789 233835 8823
rect 230397 8585 230431 8619
rect 245117 8449 245151 8483
rect 245577 8449 245611 8483
rect 247877 9537 247911 9571
rect 248245 9537 248279 9571
rect 270877 9537 270911 9571
rect 170321 8381 170355 8415
rect 266829 9469 266863 9503
rect 271061 9469 271095 9503
rect 271429 9469 271463 9503
rect 258641 9401 258675 9435
rect 267105 9401 267139 9435
rect 258917 9333 258951 9367
rect 261493 9333 261527 9367
rect 267197 9333 267231 9367
rect 270509 9333 270543 9367
rect 253305 9197 253339 9231
rect 253121 9061 253155 9095
rect 263609 9129 263643 9163
rect 258641 9061 258675 9095
rect 253305 8857 253339 8891
rect 253397 8857 253431 8891
rect 253121 8789 253155 8823
rect 253213 8789 253247 8823
rect 253213 8585 253247 8619
rect 258549 8789 258583 8823
rect 258641 8789 258675 8823
rect 261769 9061 261803 9095
rect 263701 9061 263735 9095
rect 261677 8789 261711 8823
rect 261769 8789 261803 8823
rect 258549 8585 258583 8619
rect 261769 8585 261803 8619
rect 263701 8585 263735 8619
rect 267197 8721 267231 8755
rect 268393 8789 268427 8823
rect 268393 8585 268427 8619
rect 263793 8517 263827 8551
rect 271429 8517 271463 8551
rect 253397 8449 253431 8483
rect 263609 8449 263643 8483
rect 263885 8449 263919 8483
rect 247877 8381 247911 8415
rect 272340 9537 272374 9571
rect 277869 9537 277903 9571
rect 272073 9469 272107 9503
rect 277593 9469 277627 9503
rect 273453 9333 273487 9367
rect 273729 9333 273763 9367
rect 277409 9061 277443 9095
rect 273729 8585 273763 8619
rect 277777 8585 277811 8619
rect 271521 8381 271555 8415
rect 277777 8381 277811 8415
rect 282193 9469 282227 9503
rect 278145 9265 278179 9299
rect 280813 9265 280847 9299
rect 282101 9197 282135 9231
rect 282193 9197 282227 9231
rect 282285 9469 282319 9503
rect 280997 9061 281031 9095
rect 282193 9061 282227 9095
rect 279341 8789 279375 8823
rect 279157 8721 279191 8755
rect 282193 8721 282227 8755
rect 282285 8721 282319 8755
rect 278053 8381 278087 8415
rect 282101 8381 282135 8415
rect 282193 8517 282227 8551
rect 282193 8381 282227 8415
rect 66177 8313 66211 8347
rect 203073 7837 203107 7871
rect 69112 5185 69146 5219
rect 68845 5117 68879 5151
rect 70225 4981 70259 5015
rect 225521 4437 225555 4471
rect 310989 4029 311023 4063
rect 318717 4029 318751 4063
rect 310989 3349 311023 3383
rect 312093 3349 312127 3383
rect 318717 3349 318751 3383
rect 498209 3213 498243 3247
rect 312093 3009 312127 3043
<< metal1 >>
rect 369854 617516 369860 617568
rect 369912 617556 369918 617568
rect 371142 617556 371148 617568
rect 369912 617528 371148 617556
rect 369912 617516 369918 617528
rect 371142 617516 371148 617528
rect 371200 617516 371206 617568
rect 463694 617516 463700 617568
rect 463752 617556 463758 617568
rect 464982 617556 464988 617568
rect 463752 617528 464988 617556
rect 463752 617516 463758 617528
rect 464982 617516 464988 617528
rect 465040 617516 465046 617568
rect 494054 617516 494060 617568
rect 494112 617556 494118 617568
rect 495342 617556 495348 617568
rect 494112 617528 495348 617556
rect 494112 617516 494118 617528
rect 495342 617516 495348 617528
rect 495400 617516 495406 617568
rect 3418 616836 3424 616888
rect 3476 616876 3482 616888
rect 134518 616876 134524 616888
rect 3476 616848 134524 616876
rect 3476 616836 3482 616848
rect 134518 616836 134524 616848
rect 134576 616836 134582 616888
rect 22830 616768 22836 616820
rect 22888 616808 22894 616820
rect 23382 616808 23388 616820
rect 22888 616780 23388 616808
rect 22888 616768 22894 616780
rect 23382 616768 23388 616780
rect 23440 616768 23446 616820
rect 34974 616768 34980 616820
rect 35032 616808 35038 616820
rect 35802 616808 35808 616820
rect 35032 616780 35808 616808
rect 35032 616768 35038 616780
rect 35802 616768 35808 616780
rect 35860 616768 35866 616820
rect 53006 616768 53012 616820
rect 53064 616808 53070 616820
rect 53742 616808 53748 616820
rect 53064 616780 53748 616808
rect 53064 616768 53070 616780
rect 53742 616768 53748 616780
rect 53800 616768 53806 616820
rect 77294 616768 77300 616820
rect 77352 616808 77358 616820
rect 78490 616808 78496 616820
rect 77352 616780 78496 616808
rect 77352 616768 77358 616780
rect 78490 616768 78496 616780
rect 78548 616768 78554 616820
rect 113726 616768 113732 616820
rect 113784 616808 113790 616820
rect 114370 616808 114376 616820
rect 113784 616780 114376 616808
rect 113784 616768 113790 616780
rect 114370 616768 114376 616780
rect 114428 616768 114434 616820
rect 143902 616768 143908 616820
rect 143960 616808 143966 616820
rect 299198 616808 299204 616820
rect 143960 616780 299204 616808
rect 143960 616768 143966 616780
rect 299198 616768 299204 616780
rect 299256 616768 299262 616820
rect 310606 616768 310612 616820
rect 310664 616808 310670 616820
rect 311802 616808 311808 616820
rect 310664 616780 311808 616808
rect 310664 616768 310670 616780
rect 311802 616768 311808 616780
rect 311860 616768 311866 616820
rect 313366 616768 313372 616820
rect 313424 616808 313430 616820
rect 428734 616808 428740 616820
rect 313424 616780 428740 616808
rect 313424 616768 313430 616780
rect 428734 616768 428740 616780
rect 428792 616768 428798 616820
rect 4614 616700 4620 616752
rect 4672 616740 4678 616752
rect 5442 616740 5448 616752
rect 4672 616712 5448 616740
rect 4672 616700 4678 616712
rect 5442 616700 5448 616712
rect 5500 616700 5506 616752
rect 65150 616700 65156 616752
rect 65208 616740 65214 616752
rect 66162 616740 66168 616752
rect 65208 616712 66168 616740
rect 65208 616700 65214 616712
rect 66162 616700 66168 616712
rect 66220 616700 66226 616752
rect 80422 616700 80428 616752
rect 80480 616740 80486 616752
rect 81342 616740 81348 616752
rect 80480 616712 81348 616740
rect 80480 616700 80486 616712
rect 81342 616700 81348 616712
rect 81400 616700 81406 616752
rect 114094 616700 114100 616752
rect 114152 616740 114158 616752
rect 265158 616740 265164 616752
rect 114152 616712 265164 616740
rect 114152 616700 114158 616712
rect 265158 616700 265164 616712
rect 265216 616700 265222 616752
rect 285306 616700 285312 616752
rect 285364 616740 285370 616752
rect 462038 616740 462044 616752
rect 285364 616712 462044 616740
rect 285364 616700 285370 616712
rect 462038 616700 462044 616712
rect 462096 616700 462102 616752
rect 471054 616700 471060 616752
rect 471112 616740 471118 616752
rect 471882 616740 471888 616752
rect 471112 616712 471888 616740
rect 471112 616700 471118 616712
rect 471882 616700 471888 616712
rect 471940 616700 471946 616752
rect 106734 616632 106740 616684
rect 106792 616672 106798 616684
rect 125870 616672 125876 616684
rect 106792 616644 125876 616672
rect 106792 616632 106798 616644
rect 125870 616632 125876 616644
rect 125928 616632 125934 616684
rect 131758 616632 131764 616684
rect 131816 616672 131822 616684
rect 315390 616672 315396 616684
rect 131816 616644 315396 616672
rect 131816 616632 131822 616644
rect 315390 616632 315396 616644
rect 315448 616632 315454 616684
rect 392302 616632 392308 616684
rect 392360 616672 392366 616684
rect 393222 616672 393228 616684
rect 392360 616644 393228 616672
rect 392360 616632 392366 616644
rect 393222 616632 393228 616644
rect 393280 616632 393286 616684
rect 101582 616564 101588 616616
rect 101640 616604 101646 616616
rect 322198 616604 322204 616616
rect 101640 616576 322204 616604
rect 101640 616564 101646 616576
rect 322198 616564 322204 616576
rect 322256 616564 322262 616616
rect 356054 616564 356060 616616
rect 356112 616604 356118 616616
rect 382550 616604 382556 616616
rect 356112 616576 382556 616604
rect 356112 616564 356118 616576
rect 382550 616564 382556 616576
rect 382608 616564 382614 616616
rect 36354 616496 36360 616548
rect 36412 616536 36418 616548
rect 134886 616536 134892 616548
rect 36412 616508 134892 616536
rect 36412 616496 36418 616508
rect 134886 616496 134892 616508
rect 134944 616496 134950 616548
rect 137830 616496 137836 616548
rect 137888 616536 137894 616548
rect 363598 616536 363604 616548
rect 137888 616508 363604 616536
rect 137888 616496 137894 616508
rect 363598 616496 363604 616508
rect 363656 616496 363662 616548
rect 17218 616428 17224 616480
rect 17276 616468 17282 616480
rect 128814 616468 128820 616480
rect 17276 616440 128820 616468
rect 17276 616428 17282 616440
rect 128814 616428 128820 616440
rect 128872 616428 128878 616480
rect 153838 616428 153844 616480
rect 153896 616468 153902 616480
rect 183278 616468 183284 616480
rect 153896 616440 183284 616468
rect 153896 616428 153902 616440
rect 183278 616428 183284 616440
rect 183336 616428 183342 616480
rect 184566 616428 184572 616480
rect 184624 616468 184630 616480
rect 416590 616468 416596 616480
rect 184624 616440 416596 616468
rect 184624 616428 184630 616440
rect 416590 616428 416596 616440
rect 416648 616428 416654 616480
rect 71222 616360 71228 616412
rect 71280 616400 71286 616412
rect 314102 616400 314108 616412
rect 71280 616372 314108 616400
rect 71280 616360 71286 616372
rect 314102 616360 314108 616372
rect 314160 616360 314166 616412
rect 331766 616360 331772 616412
rect 331824 616400 331830 616412
rect 371786 616400 371792 616412
rect 331824 616372 371792 616400
rect 331824 616360 331830 616372
rect 371786 616360 371792 616372
rect 371844 616360 371850 616412
rect 389818 616360 389824 616412
rect 389876 616400 389882 616412
rect 443822 616400 443828 616412
rect 389876 616372 443828 616400
rect 389876 616360 389882 616372
rect 443822 616360 443828 616372
rect 443880 616360 443886 616412
rect 110598 616292 110604 616344
rect 110656 616332 110662 616344
rect 425698 616332 425704 616344
rect 110656 616304 425704 616332
rect 110656 616292 110662 616304
rect 425698 616292 425704 616304
rect 425756 616292 425762 616344
rect 6822 616224 6828 616276
rect 6880 616264 6886 616276
rect 122742 616264 122748 616276
rect 6880 616236 122748 616264
rect 6880 616224 6886 616236
rect 122742 616224 122748 616236
rect 122800 616224 122806 616276
rect 136542 616224 136548 616276
rect 136600 616264 136606 616276
rect 452838 616264 452844 616276
rect 136600 616236 452844 616264
rect 136600 616224 136606 616236
rect 452838 616224 452844 616236
rect 452896 616224 452902 616276
rect 9858 616156 9864 616208
rect 9916 616196 9922 616208
rect 25774 616196 25780 616208
rect 9916 616168 25780 616196
rect 9916 616156 9922 616168
rect 25774 616156 25780 616168
rect 25832 616156 25838 616208
rect 28902 616156 28908 616208
rect 28960 616196 28966 616208
rect 103514 616196 103520 616208
rect 28960 616168 103520 616196
rect 28960 616156 28966 616168
rect 103514 616156 103520 616168
rect 103572 616156 103578 616208
rect 104526 616156 104532 616208
rect 104584 616196 104590 616208
rect 438302 616196 438308 616208
rect 104584 616168 438308 616196
rect 104584 616156 104590 616168
rect 438302 616156 438308 616168
rect 438360 616156 438366 616208
rect 1670 616088 1676 616140
rect 1728 616128 1734 616140
rect 359458 616128 359464 616140
rect 1728 616100 359464 616128
rect 1728 616088 1734 616100
rect 359458 616088 359464 616100
rect 359516 616088 359522 616140
rect 395338 616088 395344 616140
rect 395396 616128 395402 616140
rect 468110 616128 468116 616140
rect 395396 616100 468116 616128
rect 395396 616088 395402 616100
rect 468110 616088 468116 616100
rect 468168 616088 468174 616140
rect 78582 616020 78588 616072
rect 78640 616060 78646 616072
rect 162118 616060 162124 616072
rect 78640 616032 162124 616060
rect 78640 616020 78646 616032
rect 162118 616020 162124 616032
rect 162176 616020 162182 616072
rect 222654 616020 222660 616072
rect 222712 616060 222718 616072
rect 222712 616032 230888 616060
rect 222712 616020 222718 616032
rect 83366 615952 83372 616004
rect 83424 615992 83430 616004
rect 160738 615992 160744 616004
rect 83424 615964 160744 615992
rect 83424 615952 83430 615964
rect 160738 615952 160744 615964
rect 160796 615952 160802 616004
rect 230860 615992 230888 616032
rect 233418 616020 233424 616072
rect 233476 616060 233482 616072
rect 277302 616060 277308 616072
rect 233476 616032 277308 616060
rect 233476 616020 233482 616032
rect 277302 616020 277308 616032
rect 277360 616020 277366 616072
rect 281350 616020 281356 616072
rect 281408 616060 281414 616072
rect 404446 616060 404452 616072
rect 281408 616032 404452 616060
rect 281408 616020 281414 616032
rect 404446 616020 404452 616032
rect 404504 616020 404510 616072
rect 314010 615992 314016 616004
rect 230860 615964 314016 615992
rect 314010 615952 314016 615964
rect 314068 615952 314074 616004
rect 95510 615884 95516 615936
rect 95568 615924 95574 615936
rect 167730 615924 167736 615936
rect 95568 615896 167736 615924
rect 95568 615884 95574 615896
rect 167730 615884 167736 615896
rect 167788 615884 167794 615936
rect 262030 615884 262036 615936
rect 262088 615924 262094 615936
rect 346486 615924 346492 615936
rect 262088 615896 346492 615924
rect 262088 615884 262094 615896
rect 346486 615884 346492 615896
rect 346544 615884 346550 615936
rect 98454 615816 98460 615868
rect 98512 615856 98518 615868
rect 153194 615856 153200 615868
rect 98512 615828 153200 615856
rect 98512 615816 98518 615828
rect 153194 615816 153200 615828
rect 153252 615816 153258 615868
rect 216214 615816 216220 615868
rect 216272 615856 216278 615868
rect 289262 615856 289268 615868
rect 216272 615828 289268 615856
rect 216272 615816 216278 615828
rect 289262 615816 289268 615828
rect 289320 615816 289326 615868
rect 143810 615748 143816 615800
rect 143868 615788 143874 615800
rect 198550 615788 198556 615800
rect 143868 615760 198556 615788
rect 143868 615748 143874 615760
rect 198550 615748 198556 615760
rect 198608 615748 198614 615800
rect 210510 615748 210516 615800
rect 210568 615788 210574 615800
rect 211062 615788 211068 615800
rect 210568 615760 211068 615788
rect 210568 615748 210574 615760
rect 211062 615748 211068 615760
rect 211120 615748 211126 615800
rect 247586 615748 247592 615800
rect 247644 615788 247650 615800
rect 298462 615788 298468 615800
rect 247644 615760 298468 615788
rect 247644 615748 247650 615760
rect 298462 615748 298468 615760
rect 298520 615748 298526 615800
rect 268378 615680 268384 615732
rect 268436 615720 268442 615732
rect 313550 615720 313556 615732
rect 268436 615692 313556 615720
rect 268436 615680 268442 615692
rect 313550 615680 313556 615692
rect 313608 615680 313614 615732
rect 280246 615544 280252 615596
rect 280304 615584 280310 615596
rect 281442 615584 281448 615596
rect 280304 615556 281448 615584
rect 280304 615544 280310 615556
rect 281442 615544 281448 615556
rect 281500 615544 281506 615596
rect 334710 615544 334716 615596
rect 334768 615584 334774 615596
rect 334768 615556 335354 615584
rect 334768 615544 334774 615556
rect 335326 615516 335354 615556
rect 492950 615516 492956 615528
rect 335326 615488 492956 615516
rect 492950 615476 492956 615488
rect 493008 615476 493014 615528
rect 364242 614972 364248 614984
rect 364203 614944 364248 614972
rect 364242 614932 364248 614944
rect 364300 614932 364306 614984
rect 167549 613955 167607 613961
rect 161446 613924 167500 613952
rect 137186 613844 137192 613896
rect 137244 613884 137250 613896
rect 161446 613884 161474 613924
rect 167270 613884 167276 613896
rect 137244 613856 161474 613884
rect 167231 613856 167276 613884
rect 137244 613844 137250 613856
rect 167270 613844 167276 613856
rect 167328 613844 167334 613896
rect 167472 613893 167500 613924
rect 167549 613921 167561 613955
rect 167595 613952 167607 613955
rect 175734 613952 175740 613964
rect 167595 613924 175740 613952
rect 167595 613921 167607 613924
rect 167549 613915 167607 613921
rect 175734 613912 175740 613924
rect 175792 613912 175798 613964
rect 167457 613887 167515 613893
rect 167457 613853 167469 613887
rect 167503 613853 167515 613887
rect 167638 613884 167644 613896
rect 167599 613856 167644 613884
rect 167457 613847 167515 613853
rect 167638 613844 167644 613856
rect 167696 613844 167702 613896
rect 167733 613887 167791 613893
rect 167733 613853 167745 613887
rect 167779 613884 167791 613887
rect 167779 613856 171134 613884
rect 167779 613853 167791 613856
rect 167733 613847 167791 613853
rect 171106 613816 171134 613856
rect 175642 613816 175648 613828
rect 171106 613788 175648 613816
rect 175642 613776 175648 613788
rect 175700 613776 175706 613828
rect 167914 613748 167920 613760
rect 167875 613720 167920 613748
rect 167914 613708 167920 613720
rect 167972 613708 167978 613760
rect 182082 612756 182088 612808
rect 182140 612796 182146 612808
rect 495434 612796 495440 612808
rect 182140 612768 495440 612796
rect 182140 612756 182146 612768
rect 495434 612756 495440 612768
rect 495492 612756 495498 612808
rect 376205 611711 376263 611717
rect 376205 611677 376217 611711
rect 376251 611708 376263 611711
rect 402422 611708 402428 611720
rect 376251 611680 402428 611708
rect 376251 611677 376263 611680
rect 376205 611671 376263 611677
rect 402422 611668 402428 611680
rect 402480 611668 402486 611720
rect 237834 611532 237840 611584
rect 237892 611572 237898 611584
rect 376021 611575 376079 611581
rect 376021 611572 376033 611575
rect 237892 611544 376033 611572
rect 237892 611532 237898 611544
rect 376021 611541 376033 611544
rect 376067 611541 376079 611575
rect 376021 611535 376079 611541
rect 283392 610660 287054 610688
rect 283006 610620 283012 610632
rect 282967 610592 283012 610620
rect 283006 610580 283012 610592
rect 283064 610580 283070 610632
rect 283157 610623 283215 610629
rect 283157 610589 283169 610623
rect 283203 610620 283215 610623
rect 283392 610620 283420 610660
rect 283203 610592 283420 610620
rect 283515 610623 283573 610629
rect 283203 610589 283215 610592
rect 283157 610583 283215 610589
rect 283515 610589 283527 610623
rect 283561 610620 283573 610623
rect 284205 610623 284263 610629
rect 284205 610620 284217 610623
rect 283561 610592 284217 610620
rect 283561 610589 283573 610592
rect 283515 610583 283573 610589
rect 284205 610589 284217 610592
rect 284251 610589 284263 610623
rect 287026 610620 287054 610660
rect 435266 610620 435272 610632
rect 287026 610592 435272 610620
rect 284205 610583 284263 610589
rect 435266 610580 435272 610592
rect 435324 610580 435330 610632
rect 283282 610552 283288 610564
rect 283243 610524 283288 610552
rect 283282 610512 283288 610524
rect 283340 610512 283346 610564
rect 283374 610512 283380 610564
rect 283432 610552 283438 610564
rect 456794 610552 456800 610564
rect 283432 610524 283477 610552
rect 283576 610524 456800 610552
rect 283432 610512 283438 610524
rect 283300 610484 283328 610512
rect 283576 610484 283604 610524
rect 456794 610512 456800 610524
rect 456852 610512 456858 610564
rect 283300 610456 283604 610484
rect 283653 610487 283711 610493
rect 283653 610453 283665 610487
rect 283699 610484 283711 610487
rect 440878 610484 440884 610496
rect 283699 610456 440884 610484
rect 283699 610453 283711 610456
rect 283653 610447 283711 610453
rect 440878 610444 440884 610456
rect 440936 610444 440942 610496
rect 284205 610283 284263 610289
rect 284205 610249 284217 610283
rect 284251 610280 284263 610283
rect 434898 610280 434904 610292
rect 284251 610252 434904 610280
rect 284251 610249 284263 610252
rect 284205 610243 284263 610249
rect 434898 610240 434904 610252
rect 434956 610240 434962 610292
rect 283006 610172 283012 610224
rect 283064 610212 283070 610224
rect 419534 610212 419540 610224
rect 283064 610184 419540 610212
rect 283064 610172 283070 610184
rect 419534 610172 419540 610184
rect 419592 610172 419598 610224
rect 200853 609535 200911 609541
rect 200853 609501 200865 609535
rect 200899 609532 200911 609535
rect 386414 609532 386420 609544
rect 200899 609504 386420 609532
rect 200899 609501 200911 609504
rect 200853 609495 200911 609501
rect 386414 609492 386420 609504
rect 386472 609492 386478 609544
rect 129645 608855 129703 608861
rect 129645 608821 129657 608855
rect 129691 608852 129703 608855
rect 480254 608852 480260 608864
rect 129691 608824 480260 608852
rect 129691 608821 129703 608824
rect 129645 608815 129703 608821
rect 480254 608812 480260 608824
rect 480312 608812 480318 608864
rect 3050 608744 3056 608796
rect 3108 608784 3114 608796
rect 6178 608784 6184 608796
rect 3108 608756 6184 608784
rect 3108 608744 3114 608756
rect 6178 608744 6184 608756
rect 6236 608744 6242 608796
rect 334894 607968 334900 607980
rect 334855 607940 334900 607968
rect 334894 607928 334900 607940
rect 334952 607928 334958 607980
rect 334710 607764 334716 607776
rect 334671 607736 334716 607764
rect 334710 607724 334716 607736
rect 334768 607724 334774 607776
rect 200485 607359 200543 607365
rect 200485 607325 200497 607359
rect 200531 607356 200543 607359
rect 236454 607356 236460 607368
rect 200531 607328 236460 607356
rect 200531 607325 200543 607328
rect 200485 607319 200543 607325
rect 236454 607316 236460 607328
rect 236512 607316 236518 607368
rect 200393 607223 200451 607229
rect 200393 607189 200405 607223
rect 200439 607220 200451 607223
rect 263870 607220 263876 607232
rect 200439 607192 263876 607220
rect 200439 607189 200451 607192
rect 200393 607183 200451 607189
rect 263870 607180 263876 607192
rect 263928 607180 263934 607232
rect 228450 606889 228456 606892
rect 228444 606843 228456 606889
rect 228508 606880 228514 606892
rect 228508 606852 228544 606880
rect 228450 606840 228456 606843
rect 228508 606840 228514 606852
rect 228177 606815 228235 606821
rect 228177 606781 228189 606815
rect 228223 606781 228235 606815
rect 228177 606775 228235 606781
rect 228192 606676 228220 606775
rect 228100 606648 228220 606676
rect 229557 606679 229615 606685
rect 228100 606472 228128 606648
rect 229557 606645 229569 606679
rect 229603 606676 229615 606679
rect 310790 606676 310796 606688
rect 229603 606648 310796 606676
rect 229603 606645 229615 606648
rect 229557 606639 229615 606645
rect 310790 606636 310796 606648
rect 310848 606636 310854 606688
rect 231854 606472 231860 606484
rect 228100 606444 231860 606472
rect 231854 606432 231860 606444
rect 231912 606432 231918 606484
rect 3418 604460 3424 604512
rect 3476 604500 3482 604512
rect 55490 604500 55496 604512
rect 3476 604472 55496 604500
rect 3476 604460 3482 604472
rect 55490 604460 55496 604472
rect 55548 604460 55554 604512
rect 78490 604052 78496 604104
rect 78548 604092 78554 604104
rect 322201 604095 322259 604101
rect 322201 604092 322213 604095
rect 78548 604064 322213 604092
rect 78548 604052 78554 604064
rect 322201 604061 322213 604064
rect 322247 604061 322259 604095
rect 322201 604055 322259 604061
rect 184566 601440 184572 601452
rect 184527 601412 184572 601440
rect 184566 601400 184572 601412
rect 184624 601400 184630 601452
rect 22741 600831 22799 600837
rect 22741 600797 22753 600831
rect 22787 600828 22799 600831
rect 196434 600828 196440 600840
rect 22787 600800 196440 600828
rect 22787 600797 22799 600800
rect 22741 600791 22799 600797
rect 196434 600788 196440 600800
rect 196492 600788 196498 600840
rect 23014 600769 23020 600772
rect 23008 600723 23020 600769
rect 23072 600760 23078 600772
rect 23072 600732 23108 600760
rect 23014 600720 23020 600723
rect 23072 600720 23078 600732
rect 24121 600695 24179 600701
rect 24121 600661 24133 600695
rect 24167 600692 24179 600695
rect 142430 600692 142436 600704
rect 24167 600664 142436 600692
rect 24167 600661 24179 600664
rect 24121 600655 24179 600661
rect 142430 600652 142436 600664
rect 142488 600652 142494 600704
rect 233418 600284 233424 600296
rect 233379 600256 233424 600284
rect 233418 600244 233424 600256
rect 233476 600244 233482 600296
rect 53834 599400 53840 599412
rect 45526 599372 53840 599400
rect 3510 599292 3516 599344
rect 3568 599332 3574 599344
rect 45526 599332 45554 599372
rect 53834 599360 53840 599372
rect 53892 599360 53898 599412
rect 3568 599304 45554 599332
rect 50433 599335 50491 599341
rect 3568 599292 3574 599304
rect 50433 599301 50445 599335
rect 50479 599332 50491 599335
rect 50479 599304 55214 599332
rect 50479 599301 50491 599304
rect 50433 599295 50491 599301
rect 50336 599267 50394 599273
rect 50336 599233 50348 599267
rect 50382 599264 50394 599267
rect 50525 599267 50583 599273
rect 50382 599236 50476 599264
rect 50382 599233 50394 599236
rect 50336 599227 50394 599233
rect 50154 599060 50160 599072
rect 50115 599032 50160 599060
rect 50154 599020 50160 599032
rect 50212 599020 50218 599072
rect 50448 599060 50476 599236
rect 50525 599233 50537 599267
rect 50571 599233 50583 599267
rect 50525 599227 50583 599233
rect 50709 599267 50767 599273
rect 50709 599233 50721 599267
rect 50755 599264 50767 599267
rect 50985 599267 51043 599273
rect 50985 599264 50997 599267
rect 50755 599236 50997 599264
rect 50755 599233 50767 599236
rect 50709 599227 50767 599233
rect 50985 599233 50997 599236
rect 51031 599233 51043 599267
rect 55186 599264 55214 599304
rect 331214 599264 331220 599276
rect 55186 599236 331220 599264
rect 50985 599227 51043 599233
rect 50540 599196 50568 599227
rect 331214 599224 331220 599236
rect 331272 599224 331278 599276
rect 158898 599196 158904 599208
rect 50540 599168 158904 599196
rect 158898 599156 158904 599168
rect 158956 599156 158962 599208
rect 50985 599131 51043 599137
rect 50985 599097 50997 599131
rect 51031 599128 51043 599131
rect 158990 599128 158996 599140
rect 51031 599100 158996 599128
rect 51031 599097 51043 599100
rect 50985 599091 51043 599097
rect 158990 599088 158996 599100
rect 159048 599128 159054 599140
rect 159048 599100 161474 599128
rect 159048 599088 159054 599100
rect 79226 599060 79232 599072
rect 50448 599032 79232 599060
rect 79226 599020 79232 599032
rect 79284 599020 79290 599072
rect 161446 599060 161474 599100
rect 325602 599060 325608 599072
rect 161446 599032 325608 599060
rect 325602 599020 325608 599032
rect 325660 599020 325666 599072
rect 314194 598952 314200 599004
rect 314252 598992 314258 599004
rect 495434 598992 495440 599004
rect 314252 598964 495440 598992
rect 314252 598952 314258 598964
rect 495434 598952 495440 598964
rect 495492 598952 495498 599004
rect 247586 596680 247592 596692
rect 247547 596652 247592 596680
rect 247586 596640 247592 596652
rect 247644 596640 247650 596692
rect 206002 596544 206008 596556
rect 205963 596516 206008 596544
rect 206002 596504 206008 596516
rect 206060 596504 206066 596556
rect 205450 596340 205456 596352
rect 205411 596312 205456 596340
rect 205450 596300 205456 596312
rect 205508 596300 205514 596352
rect 205818 596340 205824 596352
rect 205779 596312 205824 596340
rect 205818 596300 205824 596312
rect 205876 596300 205882 596352
rect 205910 596300 205916 596352
rect 205968 596340 205974 596352
rect 205968 596312 206013 596340
rect 205968 596300 205974 596312
rect 2774 595008 2780 595060
rect 2832 595048 2838 595060
rect 5166 595048 5172 595060
rect 2832 595020 5172 595048
rect 2832 595008 2838 595020
rect 5166 595008 5172 595020
rect 5224 595008 5230 595060
rect 492950 591240 492956 591252
rect 492911 591212 492956 591240
rect 492950 591200 492956 591212
rect 493008 591200 493014 591252
rect 494330 591036 494336 591048
rect 494291 591008 494336 591036
rect 494330 590996 494336 591008
rect 494388 590996 494394 591048
rect 111886 590928 111892 590980
rect 111944 590968 111950 590980
rect 494066 590971 494124 590977
rect 494066 590968 494078 590971
rect 111944 590940 494078 590968
rect 111944 590928 111950 590940
rect 494066 590937 494078 590940
rect 494112 590937 494124 590971
rect 494066 590931 494124 590937
rect 419534 590628 419540 590640
rect 419495 590600 419540 590628
rect 419534 590588 419540 590600
rect 419592 590628 419598 590640
rect 419592 590600 422294 590628
rect 419592 590588 419598 590600
rect 419350 590560 419356 590572
rect 419311 590532 419356 590560
rect 419350 590520 419356 590532
rect 419408 590520 419414 590572
rect 422266 590560 422294 590600
rect 435358 590560 435364 590572
rect 422266 590532 435364 590560
rect 435358 590520 435364 590532
rect 435416 590520 435422 590572
rect 419626 590356 419632 590368
rect 419587 590328 419632 590356
rect 419626 590316 419632 590328
rect 419684 590316 419690 590368
rect 463436 587336 470594 587364
rect 463436 587308 463464 587336
rect 463418 587296 463424 587308
rect 463331 587268 463424 587296
rect 463418 587256 463424 587268
rect 463476 587256 463482 587308
rect 463510 587256 463516 587308
rect 463568 587296 463574 587308
rect 470566 587296 470594 587336
rect 495526 587296 495532 587308
rect 463568 587268 463613 587296
rect 470566 587268 495532 587296
rect 463568 587256 463574 587268
rect 495526 587256 495532 587268
rect 495584 587256 495590 587308
rect 463142 587228 463148 587240
rect 463103 587200 463148 587228
rect 463142 587188 463148 587200
rect 463200 587188 463206 587240
rect 203978 587052 203984 587104
rect 204036 587092 204042 587104
rect 463237 587095 463295 587101
rect 463237 587092 463249 587095
rect 204036 587064 463249 587092
rect 204036 587052 204042 587064
rect 463237 587061 463249 587064
rect 463283 587061 463295 587095
rect 463237 587055 463295 587061
rect 463697 587095 463755 587101
rect 463697 587061 463709 587095
rect 463743 587092 463755 587095
rect 463743 587064 463924 587092
rect 463743 587061 463755 587064
rect 463697 587055 463755 587061
rect 416682 586848 416688 586900
rect 416740 586888 416746 586900
rect 463896 586888 463924 587064
rect 416740 586860 463924 586888
rect 416740 586848 416746 586860
rect 2774 586508 2780 586560
rect 2832 586548 2838 586560
rect 4890 586548 4896 586560
rect 2832 586520 4896 586548
rect 2832 586508 2838 586520
rect 4890 586508 4896 586520
rect 4948 586508 4954 586560
rect 313366 586208 313372 586220
rect 313327 586180 313372 586208
rect 313366 586168 313372 586180
rect 313424 586168 313430 586220
rect 4798 585556 4804 585608
rect 4856 585596 4862 585608
rect 410337 585599 410395 585605
rect 410337 585596 410349 585599
rect 4856 585568 410349 585596
rect 4856 585556 4862 585568
rect 410337 585565 410349 585568
rect 410383 585565 410395 585599
rect 410337 585559 410395 585565
rect 106734 584712 106740 584724
rect 106695 584684 106740 584712
rect 106734 584672 106740 584684
rect 106792 584672 106798 584724
rect 206002 584400 206008 584452
rect 206060 584440 206066 584452
rect 262490 584440 262496 584452
rect 206060 584412 262496 584440
rect 206060 584400 206066 584412
rect 262490 584400 262496 584412
rect 262548 584400 262554 584452
rect 142062 583992 142068 584044
rect 142120 584032 142126 584044
rect 201589 584035 201647 584041
rect 201589 584032 201601 584035
rect 142120 584004 201601 584032
rect 142120 583992 142126 584004
rect 201589 584001 201601 584004
rect 201635 584001 201647 584035
rect 201589 583995 201647 584001
rect 201313 583967 201371 583973
rect 201313 583933 201325 583967
rect 201359 583933 201371 583967
rect 201494 583964 201500 583976
rect 201455 583936 201500 583964
rect 201313 583927 201371 583933
rect 201328 583896 201356 583927
rect 201494 583924 201500 583936
rect 201552 583924 201558 583976
rect 206002 583896 206008 583908
rect 201328 583868 206008 583896
rect 206002 583856 206008 583868
rect 206060 583856 206066 583908
rect 201954 583828 201960 583840
rect 201915 583800 201960 583828
rect 201954 583788 201960 583800
rect 202012 583788 202018 583840
rect 405918 583420 405924 583432
rect 405879 583392 405924 583420
rect 405918 583380 405924 583392
rect 405976 583380 405982 583432
rect 28902 580728 28908 580780
rect 28960 580768 28966 580780
rect 482557 580771 482615 580777
rect 482557 580768 482569 580771
rect 28960 580740 482569 580768
rect 28960 580728 28966 580740
rect 482557 580737 482569 580740
rect 482603 580737 482615 580771
rect 482557 580731 482615 580737
rect 482646 580700 482652 580712
rect 482607 580672 482652 580700
rect 482646 580660 482652 580672
rect 482704 580660 482710 580712
rect 482738 580660 482744 580712
rect 482796 580700 482802 580712
rect 482796 580672 482841 580700
rect 482796 580660 482802 580672
rect 372706 580524 372712 580576
rect 372764 580564 372770 580576
rect 482189 580567 482247 580573
rect 482189 580564 482201 580567
rect 372764 580536 482201 580564
rect 372764 580524 372770 580536
rect 482189 580533 482201 580536
rect 482235 580533 482247 580567
rect 482189 580527 482247 580533
rect 396905 579139 396963 579145
rect 396905 579105 396917 579139
rect 396951 579136 396963 579139
rect 396951 579108 402974 579136
rect 396951 579105 396963 579108
rect 396905 579099 396963 579105
rect 113637 579071 113695 579077
rect 113637 579037 113649 579071
rect 113683 579068 113695 579071
rect 291194 579068 291200 579080
rect 113683 579040 291200 579068
rect 113683 579037 113695 579040
rect 113637 579031 113695 579037
rect 291194 579028 291200 579040
rect 291252 579028 291258 579080
rect 396629 579003 396687 579009
rect 396629 579000 396641 579003
rect 393286 578972 396641 579000
rect 121362 578892 121368 578944
rect 121420 578932 121426 578944
rect 393286 578932 393314 578972
rect 396629 578969 396641 578972
rect 396675 578969 396687 579003
rect 396629 578963 396687 578969
rect 396261 578935 396319 578941
rect 396261 578932 396273 578935
rect 121420 578904 393314 578932
rect 394804 578904 396273 578932
rect 121420 578892 121426 578904
rect 180426 578688 180432 578740
rect 180484 578728 180490 578740
rect 394804 578728 394832 578904
rect 396261 578901 396273 578904
rect 396307 578901 396319 578935
rect 396261 578895 396319 578901
rect 396718 578892 396724 578944
rect 396776 578932 396782 578944
rect 402946 578932 402974 579108
rect 403434 578932 403440 578944
rect 396776 578904 396821 578932
rect 402946 578904 403440 578932
rect 396776 578892 396782 578904
rect 403434 578892 403440 578904
rect 403492 578932 403498 578944
rect 482738 578932 482744 578944
rect 403492 578904 482744 578932
rect 403492 578892 403498 578904
rect 482738 578892 482744 578904
rect 482796 578892 482802 578944
rect 180484 578700 394832 578728
rect 180484 578688 180490 578700
rect 3602 578348 3608 578400
rect 3660 578388 3666 578400
rect 248233 578391 248291 578397
rect 248233 578388 248245 578391
rect 3660 578360 248245 578388
rect 3660 578348 3666 578360
rect 248233 578357 248245 578360
rect 248279 578357 248291 578391
rect 248233 578351 248291 578357
rect 2774 577260 2780 577312
rect 2832 577300 2838 577312
rect 4982 577300 4988 577312
rect 2832 577272 4988 577300
rect 2832 577260 2838 577272
rect 4982 577260 4988 577272
rect 5040 577260 5046 577312
rect 247678 576920 247684 576972
rect 247736 576960 247742 576972
rect 423769 576963 423827 576969
rect 423769 576960 423781 576963
rect 247736 576932 423781 576960
rect 247736 576920 247742 576932
rect 423769 576929 423781 576932
rect 423815 576929 423827 576963
rect 423769 576923 423827 576929
rect 233326 576852 233332 576904
rect 233384 576892 233390 576904
rect 423401 576895 423459 576901
rect 423401 576892 423413 576895
rect 233384 576864 423413 576892
rect 233384 576852 233390 576864
rect 423401 576861 423413 576864
rect 423447 576861 423459 576895
rect 423582 576892 423588 576904
rect 423543 576864 423588 576892
rect 423401 576855 423459 576861
rect 423582 576852 423588 576864
rect 423640 576852 423646 576904
rect 66162 576172 66168 576224
rect 66220 576212 66226 576224
rect 417513 576215 417571 576221
rect 417513 576212 417525 576215
rect 66220 576184 417525 576212
rect 66220 576172 66226 576184
rect 417513 576181 417525 576184
rect 417559 576181 417571 576215
rect 417513 576175 417571 576181
rect 43070 572704 43076 572756
rect 43128 572744 43134 572756
rect 495434 572744 495440 572756
rect 43128 572716 495440 572744
rect 43128 572704 43134 572716
rect 495434 572704 495440 572716
rect 495492 572704 495498 572756
rect 231854 572132 231860 572144
rect 196452 572104 231860 572132
rect 196452 572076 196480 572104
rect 231854 572092 231860 572104
rect 231912 572092 231918 572144
rect 196434 572064 196440 572076
rect 196395 572036 196440 572064
rect 196434 572024 196440 572036
rect 196492 572024 196498 572076
rect 196704 572067 196762 572073
rect 196704 572033 196716 572067
rect 196750 572064 196762 572067
rect 422938 572064 422944 572076
rect 196750 572036 422944 572064
rect 196750 572033 196762 572036
rect 196704 572027 196762 572033
rect 422938 572024 422944 572036
rect 422996 572024 423002 572076
rect 369397 571999 369455 572005
rect 369397 571996 369409 571999
rect 354646 571968 369409 571996
rect 213822 571888 213828 571940
rect 213880 571928 213886 571940
rect 354646 571928 354674 571968
rect 369397 571965 369409 571968
rect 369443 571965 369455 571999
rect 369397 571959 369455 571965
rect 213880 571900 354674 571928
rect 369136 571900 373994 571928
rect 213880 571888 213886 571900
rect 197817 571863 197875 571869
rect 197817 571829 197829 571863
rect 197863 571860 197875 571863
rect 369136 571860 369164 571900
rect 197863 571832 369164 571860
rect 373966 571860 373994 571900
rect 445662 571860 445668 571872
rect 373966 571832 445668 571860
rect 197863 571829 197875 571832
rect 197817 571823 197875 571829
rect 445662 571820 445668 571832
rect 445720 571820 445726 571872
rect 236454 571112 236460 571124
rect 236415 571084 236460 571112
rect 236454 571072 236460 571084
rect 236512 571072 236518 571124
rect 237558 570976 237564 570988
rect 237616 570985 237622 570988
rect 237528 570948 237564 570976
rect 237558 570936 237564 570948
rect 237616 570939 237628 570985
rect 237834 570976 237840 570988
rect 237795 570948 237840 570976
rect 237616 570936 237622 570939
rect 237834 570936 237840 570948
rect 237892 570936 237898 570988
rect 285306 570976 285312 570988
rect 285267 570948 285312 570976
rect 285306 570936 285312 570948
rect 285364 570936 285370 570988
rect 236454 570732 236460 570784
rect 236512 570772 236518 570784
rect 417878 570772 417884 570784
rect 236512 570744 417884 570772
rect 236512 570732 236518 570744
rect 417878 570732 417884 570744
rect 417936 570732 417942 570784
rect 376478 569276 376484 569288
rect 376439 569248 376484 569276
rect 376478 569236 376484 569248
rect 376536 569236 376542 569288
rect 473722 567100 473728 567112
rect 473683 567072 473728 567100
rect 473722 567060 473728 567072
rect 473780 567060 473786 567112
rect 473906 567100 473912 567112
rect 473867 567072 473912 567100
rect 473906 567060 473912 567072
rect 473964 567060 473970 567112
rect 451918 566924 451924 566976
rect 451976 566964 451982 566976
rect 473817 566967 473875 566973
rect 473817 566964 473829 566967
rect 451976 566936 473829 566964
rect 451976 566924 451982 566936
rect 473817 566933 473829 566936
rect 473863 566933 473875 566967
rect 473817 566927 473875 566933
rect 78582 566216 78588 566228
rect 78543 566188 78588 566216
rect 78582 566176 78588 566188
rect 78640 566176 78646 566228
rect 80977 566083 81035 566089
rect 80977 566080 80989 566083
rect 75656 566052 80989 566080
rect 75656 566021 75684 566052
rect 80977 566049 80989 566052
rect 81023 566049 81035 566083
rect 80977 566043 81035 566049
rect 75641 566015 75699 566021
rect 75641 565981 75653 566015
rect 75687 565981 75699 566015
rect 75641 565975 75699 565981
rect 75825 566015 75883 566021
rect 75825 565981 75837 566015
rect 75871 565981 75883 566015
rect 76010 566015 76068 566021
rect 75825 565975 75883 565981
rect 75918 565993 75976 565999
rect 75840 565876 75868 565975
rect 75918 565959 75930 565993
rect 75964 565959 75976 565993
rect 76010 565981 76022 566015
rect 76056 566012 76068 566015
rect 233694 566012 233700 566024
rect 76056 565984 233700 566012
rect 76056 565981 76068 565984
rect 76010 565975 76068 565981
rect 233694 565972 233700 565984
rect 233752 565972 233758 566024
rect 325602 566012 325608 566024
rect 325563 565984 325608 566012
rect 325602 565972 325608 565984
rect 325660 565972 325666 566024
rect 325786 566012 325792 566024
rect 325747 565984 325792 566012
rect 325786 565972 325792 565984
rect 325844 565972 325850 566024
rect 75918 565956 75976 565959
rect 75914 565904 75920 565956
rect 75972 565904 75978 565956
rect 76282 565944 76288 565956
rect 76243 565916 76288 565944
rect 76282 565904 76288 565916
rect 76340 565904 76346 565956
rect 208302 565944 208308 565956
rect 80900 565916 208308 565944
rect 80900 565876 80928 565916
rect 208302 565904 208308 565916
rect 208360 565904 208366 565956
rect 325510 565944 325516 565956
rect 325471 565916 325516 565944
rect 325510 565904 325516 565916
rect 325568 565904 325574 565956
rect 75840 565848 80928 565876
rect 80977 565879 81035 565885
rect 80977 565845 80989 565879
rect 81023 565876 81035 565879
rect 158438 565876 158444 565888
rect 81023 565848 158444 565876
rect 81023 565845 81035 565848
rect 80977 565839 81035 565845
rect 158438 565836 158444 565848
rect 158496 565836 158502 565888
rect 15010 561728 15016 561740
rect 14971 561700 15016 561728
rect 15010 561688 15016 561700
rect 15068 561688 15074 561740
rect 15473 561731 15531 561737
rect 15473 561697 15485 561731
rect 15519 561728 15531 561731
rect 51442 561728 51448 561740
rect 15519 561700 51448 561728
rect 15519 561697 15531 561700
rect 15473 561691 15531 561697
rect 51442 561688 51448 561700
rect 51500 561688 51506 561740
rect 15197 561663 15255 561669
rect 15197 561629 15209 561663
rect 15243 561629 15255 561663
rect 15197 561623 15255 561629
rect 15212 561524 15240 561623
rect 15286 561620 15292 561672
rect 15344 561660 15350 561672
rect 15565 561663 15623 561669
rect 15344 561632 15389 561660
rect 15344 561620 15350 561632
rect 15565 561629 15577 561663
rect 15611 561629 15623 561663
rect 15565 561623 15623 561629
rect 16117 561663 16175 561669
rect 16117 561629 16129 561663
rect 16163 561660 16175 561663
rect 258902 561660 258908 561672
rect 16163 561632 258908 561660
rect 16163 561629 16175 561632
rect 16117 561623 16175 561629
rect 15580 561592 15608 561623
rect 258902 561620 258908 561632
rect 258960 561620 258966 561672
rect 123386 561592 123392 561604
rect 15580 561564 123392 561592
rect 123386 561552 123392 561564
rect 123444 561552 123450 561604
rect 16117 561527 16175 561533
rect 16117 561524 16129 561527
rect 15212 561496 16129 561524
rect 16117 561493 16129 561496
rect 16163 561493 16175 561527
rect 16117 561487 16175 561493
rect 203978 559144 203984 559156
rect 203939 559116 203984 559144
rect 203978 559104 203984 559116
rect 204036 559104 204042 559156
rect 204165 559011 204223 559017
rect 204165 558977 204177 559011
rect 204211 559008 204223 559011
rect 255682 559008 255688 559020
rect 204211 558980 255688 559008
rect 204211 558977 204223 558980
rect 204165 558971 204223 558977
rect 255682 558968 255688 558980
rect 255740 558968 255746 559020
rect 2866 558900 2872 558952
rect 2924 558940 2930 558952
rect 101398 558940 101404 558952
rect 2924 558912 101404 558940
rect 2924 558900 2930 558912
rect 101398 558900 101404 558912
rect 101456 558900 101462 558952
rect 204346 558940 204352 558952
rect 204307 558912 204352 558940
rect 204346 558900 204352 558912
rect 204404 558900 204410 558952
rect 403434 557376 403440 557388
rect 403395 557348 403440 557376
rect 403434 557336 403440 557348
rect 403492 557336 403498 557388
rect 403253 557243 403311 557249
rect 403253 557240 403265 557243
rect 393286 557212 403265 557240
rect 82722 557132 82728 557184
rect 82780 557172 82786 557184
rect 393286 557172 393314 557212
rect 403253 557209 403265 557212
rect 403299 557209 403311 557243
rect 403253 557203 403311 557209
rect 402885 557175 402943 557181
rect 402885 557172 402897 557175
rect 82780 557144 393314 557172
rect 398116 557144 402897 557172
rect 82780 557132 82786 557144
rect 327258 556928 327264 556980
rect 327316 556968 327322 556980
rect 398116 556968 398144 557144
rect 402885 557141 402897 557144
rect 402931 557141 402943 557175
rect 402885 557135 402943 557141
rect 403342 557132 403348 557184
rect 403400 557172 403406 557184
rect 403400 557144 403445 557172
rect 403400 557132 403406 557144
rect 327316 556940 398144 556968
rect 327316 556928 327322 556940
rect 169956 556872 171134 556900
rect 169956 556841 169984 556872
rect 169941 556835 169999 556841
rect 169941 556801 169953 556835
rect 169987 556801 169999 556835
rect 169941 556795 169999 556801
rect 170125 556835 170183 556841
rect 170125 556801 170137 556835
rect 170171 556801 170183 556835
rect 171106 556832 171134 556872
rect 331490 556832 331496 556844
rect 171106 556804 331496 556832
rect 170125 556795 170183 556801
rect 170140 556764 170168 556795
rect 331490 556792 331496 556804
rect 331548 556792 331554 556844
rect 310606 556764 310612 556776
rect 170140 556736 310612 556764
rect 310606 556724 310612 556736
rect 310664 556724 310670 556776
rect 169849 556699 169907 556705
rect 169849 556665 169861 556699
rect 169895 556696 169907 556699
rect 316678 556696 316684 556708
rect 169895 556668 316684 556696
rect 169895 556665 169907 556668
rect 169849 556659 169907 556665
rect 316678 556656 316684 556668
rect 316736 556656 316742 556708
rect 403434 556180 403440 556232
rect 403492 556220 403498 556232
rect 406010 556220 406016 556232
rect 403492 556192 406016 556220
rect 403492 556180 403498 556192
rect 406010 556180 406016 556192
rect 406068 556180 406074 556232
rect 304905 555135 304963 555141
rect 304905 555101 304917 555135
rect 304951 555132 304963 555135
rect 313918 555132 313924 555144
rect 304951 555104 313924 555132
rect 304951 555101 304963 555104
rect 304905 555095 304963 555101
rect 313918 555092 313924 555104
rect 313976 555092 313982 555144
rect 2774 554752 2780 554804
rect 2832 554792 2838 554804
rect 6270 554792 6276 554804
rect 2832 554764 6276 554792
rect 2832 554752 2838 554764
rect 6270 554752 6276 554764
rect 6328 554752 6334 554804
rect 316770 554752 316776 554804
rect 316828 554792 316834 554804
rect 495434 554792 495440 554804
rect 316828 554764 495440 554792
rect 316828 554752 316834 554764
rect 495434 554752 495440 554764
rect 495492 554752 495498 554804
rect 330846 554044 330852 554056
rect 330807 554016 330852 554044
rect 330846 554004 330852 554016
rect 330904 554004 330910 554056
rect 268286 553528 268292 553580
rect 268344 553577 268350 553580
rect 268344 553571 268393 553577
rect 268344 553537 268347 553571
rect 268381 553537 268393 553571
rect 268344 553531 268393 553537
rect 268473 553571 268531 553577
rect 268473 553537 268485 553571
rect 268519 553537 268531 553571
rect 268473 553531 268531 553537
rect 268344 553528 268350 553531
rect 268488 553500 268516 553531
rect 268562 553528 268568 553580
rect 268620 553568 268626 553580
rect 268746 553568 268752 553580
rect 268620 553540 268665 553568
rect 268707 553540 268752 553568
rect 268620 553528 268626 553540
rect 268746 553528 268752 553540
rect 268804 553528 268810 553580
rect 268838 553528 268844 553580
rect 268896 553568 268902 553580
rect 268896 553540 268941 553568
rect 268896 553528 268902 553540
rect 447778 553500 447784 553512
rect 268488 553472 447784 553500
rect 447778 553460 447784 553472
rect 447836 553460 447842 553512
rect 268197 553435 268255 553441
rect 268197 553401 268209 553435
rect 268243 553432 268255 553435
rect 376202 553432 376208 553444
rect 268243 553404 376208 553432
rect 268243 553401 268255 553404
rect 268197 553395 268255 553401
rect 376202 553392 376208 553404
rect 376260 553392 376266 553444
rect 434898 551877 434904 551880
rect 434896 551868 434904 551877
rect 434859 551840 434904 551868
rect 434896 551831 434904 551840
rect 434898 551828 434904 551831
rect 434956 551828 434962 551880
rect 435266 551868 435272 551880
rect 435227 551840 435272 551868
rect 435266 551828 435272 551840
rect 435324 551828 435330 551880
rect 435358 551828 435364 551880
rect 435416 551868 435422 551880
rect 435416 551840 435461 551868
rect 435416 551828 435422 551840
rect 434990 551800 434996 551812
rect 434951 551772 434996 551800
rect 434990 551760 434996 551772
rect 435048 551760 435054 551812
rect 435082 551760 435088 551812
rect 435140 551800 435146 551812
rect 435140 551772 435185 551800
rect 435140 551760 435146 551772
rect 434714 551732 434720 551744
rect 434675 551704 434720 551732
rect 434714 551692 434720 551704
rect 434772 551692 434778 551744
rect 311158 549244 311164 549296
rect 311216 549284 311222 549296
rect 495434 549284 495440 549296
rect 311216 549256 495440 549284
rect 311216 549244 311222 549256
rect 495434 549244 495440 549256
rect 495492 549244 495498 549296
rect 231854 548672 231860 548684
rect 231815 548644 231860 548672
rect 231854 548632 231860 548644
rect 231912 548632 231918 548684
rect 231872 548604 231900 548632
rect 260650 548604 260656 548616
rect 231872 548576 260656 548604
rect 260650 548564 260656 548576
rect 260708 548564 260714 548616
rect 232130 548545 232136 548548
rect 232124 548499 232136 548545
rect 232188 548536 232194 548548
rect 279234 548536 279240 548548
rect 232188 548508 232224 548536
rect 277366 548508 279240 548536
rect 232130 548496 232136 548499
rect 232188 548496 232194 548508
rect 233237 548471 233295 548477
rect 233237 548437 233249 548471
rect 233283 548468 233295 548471
rect 277366 548468 277394 548508
rect 279234 548496 279240 548508
rect 279292 548536 279298 548548
rect 343634 548536 343640 548548
rect 279292 548508 343640 548536
rect 279292 548496 279298 548508
rect 343634 548496 343640 548508
rect 343692 548496 343698 548548
rect 233283 548440 277394 548468
rect 233283 548437 233295 548440
rect 233237 548431 233295 548437
rect 380618 547516 380624 547528
rect 380579 547488 380624 547516
rect 380618 547476 380624 547488
rect 380676 547476 380682 547528
rect 119522 547408 119528 547460
rect 119580 547448 119586 547460
rect 380354 547451 380412 547457
rect 380354 547448 380366 547451
rect 119580 547420 380366 547448
rect 119580 547408 119586 547420
rect 380354 547417 380366 547420
rect 380400 547417 380412 547451
rect 380354 547411 380412 547417
rect 379238 547380 379244 547392
rect 379199 547352 379244 547380
rect 379238 547340 379244 547352
rect 379296 547340 379302 547392
rect 121822 546836 121828 546848
rect 121783 546808 121828 546836
rect 121822 546796 121828 546808
rect 121880 546796 121886 546848
rect 3142 545096 3148 545148
rect 3200 545136 3206 545148
rect 265066 545136 265072 545148
rect 3200 545108 265072 545136
rect 3200 545096 3206 545108
rect 265066 545096 265072 545108
rect 265124 545096 265130 545148
rect 363506 545096 363512 545148
rect 363564 545136 363570 545148
rect 495434 545136 495440 545148
rect 363564 545108 495440 545136
rect 363564 545096 363570 545108
rect 495434 545096 495440 545108
rect 495492 545096 495498 545148
rect 412606 544292 422294 544320
rect 3418 544212 3424 544264
rect 3476 544252 3482 544264
rect 412606 544252 412634 544292
rect 416590 544252 416596 544264
rect 3476 544224 412634 544252
rect 416551 544224 416596 544252
rect 3476 544212 3482 544224
rect 416590 544212 416596 544224
rect 416648 544212 416654 544264
rect 422266 544252 422294 544292
rect 445021 544255 445079 544261
rect 445021 544252 445033 544255
rect 422266 544224 445033 544252
rect 445021 544221 445033 544224
rect 445067 544221 445079 544255
rect 445021 544215 445079 544221
rect 334710 543844 334716 543856
rect 157444 543816 334716 543844
rect 157444 543788 157472 543816
rect 334710 543804 334716 543816
rect 334768 543804 334774 543856
rect 157242 543776 157248 543788
rect 157203 543748 157248 543776
rect 157242 543736 157248 543748
rect 157300 543736 157306 543788
rect 157426 543776 157432 543788
rect 157387 543748 157432 543776
rect 157426 543736 157432 543748
rect 157484 543736 157490 543788
rect 157518 543736 157524 543788
rect 157576 543776 157582 543788
rect 157613 543779 157671 543785
rect 157613 543776 157625 543779
rect 157576 543748 157625 543776
rect 157576 543736 157582 543748
rect 157613 543745 157625 543748
rect 157659 543745 157671 543779
rect 469582 543776 469588 543788
rect 157613 543739 157671 543745
rect 157720 543748 469588 543776
rect 157260 543708 157288 543736
rect 157720 543708 157748 543748
rect 469582 543736 469588 543748
rect 469640 543736 469646 543788
rect 157260 543680 157748 543708
rect 330846 542308 330852 542360
rect 330904 542348 330910 542360
rect 495434 542348 495440 542360
rect 330904 542320 495440 542348
rect 330904 542308 330910 542320
rect 495434 542308 495440 542320
rect 495492 542308 495498 542360
rect 119522 541736 119528 541748
rect 119483 541708 119528 541736
rect 119522 541696 119528 541708
rect 119580 541696 119586 541748
rect 123294 541668 123300 541680
rect 119724 541640 123300 541668
rect 119724 541609 119752 541640
rect 123294 541628 123300 541640
rect 123352 541668 123358 541680
rect 123352 541640 132494 541668
rect 123352 541628 123358 541640
rect 119709 541603 119767 541609
rect 119709 541569 119721 541603
rect 119755 541569 119767 541603
rect 119709 541563 119767 541569
rect 119801 541603 119859 541609
rect 119801 541569 119813 541603
rect 119847 541600 119859 541603
rect 132466 541600 132494 541640
rect 379238 541600 379244 541612
rect 119847 541572 122834 541600
rect 132466 541572 379244 541600
rect 119847 541569 119859 541572
rect 119801 541563 119859 541569
rect 120074 541532 120080 541544
rect 120035 541504 120080 541532
rect 120074 541492 120080 541504
rect 120132 541492 120138 541544
rect 122806 541532 122834 541572
rect 379238 541560 379244 541572
rect 379296 541560 379302 541612
rect 367738 541532 367744 541544
rect 122806 541504 367744 541532
rect 367738 541492 367744 541504
rect 367796 541492 367802 541544
rect 119982 541464 119988 541476
rect 119943 541436 119988 541464
rect 119982 541424 119988 541436
rect 120040 541424 120046 541476
rect 2866 540948 2872 541000
rect 2924 540988 2930 541000
rect 388438 540988 388444 541000
rect 2924 540960 388444 540988
rect 2924 540948 2930 540960
rect 388438 540948 388444 540960
rect 388496 540948 388502 541000
rect 158456 540552 161474 540580
rect 158456 540524 158484 540552
rect 158438 540512 158444 540524
rect 158399 540484 158444 540512
rect 158438 540472 158444 540484
rect 158496 540472 158502 540524
rect 158622 540512 158628 540524
rect 158583 540484 158628 540512
rect 158622 540472 158628 540484
rect 158680 540472 158686 540524
rect 158717 540515 158775 540521
rect 158717 540481 158729 540515
rect 158763 540481 158775 540515
rect 158717 540475 158775 540481
rect 158810 540505 158868 540511
rect 158732 540388 158760 540475
rect 158810 540471 158822 540505
rect 158856 540471 158868 540505
rect 158810 540465 158868 540471
rect 158824 540388 158852 540465
rect 161446 540444 161474 540552
rect 221458 540444 221464 540456
rect 161446 540416 221464 540444
rect 221458 540404 221464 540416
rect 221516 540404 221522 540456
rect 158714 540336 158720 540388
rect 158772 540336 158778 540388
rect 158806 540336 158812 540388
rect 158864 540336 158870 540388
rect 159082 540376 159088 540388
rect 159043 540348 159088 540376
rect 159082 540336 159088 540348
rect 159140 540336 159146 540388
rect 158622 540268 158628 540320
rect 158680 540308 158686 540320
rect 273898 540308 273904 540320
rect 158680 540280 273904 540308
rect 158680 540268 158686 540280
rect 273898 540268 273904 540280
rect 273956 540268 273962 540320
rect 462314 539520 462320 539572
rect 462372 539560 462378 539572
rect 463142 539560 463148 539572
rect 462372 539532 463148 539560
rect 462372 539520 462378 539532
rect 463142 539520 463148 539532
rect 463200 539520 463206 539572
rect 59357 539427 59415 539433
rect 59357 539393 59369 539427
rect 59403 539393 59415 539427
rect 59357 539387 59415 539393
rect 59372 539288 59400 539387
rect 59446 539384 59452 539436
rect 59504 539424 59510 539436
rect 463418 539424 463424 539436
rect 59504 539396 463424 539424
rect 59504 539384 59510 539396
rect 463418 539384 463424 539396
rect 463476 539384 463482 539436
rect 59725 539359 59783 539365
rect 59725 539325 59737 539359
rect 59771 539356 59783 539359
rect 462314 539356 462320 539368
rect 59771 539328 462320 539356
rect 59771 539325 59783 539328
rect 59725 539319 59783 539325
rect 462314 539316 462320 539328
rect 462372 539316 462378 539368
rect 326338 539288 326344 539300
rect 59372 539260 326344 539288
rect 326338 539248 326344 539260
rect 326396 539248 326402 539300
rect 59170 539220 59176 539232
rect 59131 539192 59176 539220
rect 59170 539180 59176 539192
rect 59228 539180 59234 539232
rect 59630 539220 59636 539232
rect 59591 539192 59636 539220
rect 59630 539180 59636 539192
rect 59688 539180 59694 539232
rect 6362 537684 6368 537736
rect 6420 537724 6426 537736
rect 17313 537727 17371 537733
rect 17313 537724 17325 537727
rect 6420 537696 17325 537724
rect 6420 537684 6426 537696
rect 17313 537693 17325 537696
rect 17359 537693 17371 537727
rect 17313 537687 17371 537693
rect 229002 537684 229008 537736
rect 229060 537724 229066 537736
rect 441893 537727 441951 537733
rect 441893 537724 441905 537727
rect 229060 537696 441905 537724
rect 229060 537684 229066 537696
rect 441893 537693 441905 537696
rect 441939 537693 441951 537727
rect 441893 537687 441951 537693
rect 3142 536800 3148 536852
rect 3200 536840 3206 536852
rect 6730 536840 6736 536852
rect 3200 536812 6736 536840
rect 3200 536800 3206 536812
rect 6730 536800 6736 536812
rect 6788 536800 6794 536852
rect 176930 536800 176936 536852
rect 176988 536840 176994 536852
rect 495434 536840 495440 536852
rect 176988 536812 495440 536840
rect 176988 536800 176994 536812
rect 495434 536800 495440 536812
rect 495492 536800 495498 536852
rect 3510 536596 3516 536648
rect 3568 536636 3574 536648
rect 327905 536639 327963 536645
rect 327905 536636 327917 536639
rect 3568 536608 327917 536636
rect 3568 536596 3574 536608
rect 327905 536605 327917 536608
rect 327951 536605 327963 536639
rect 327905 536599 327963 536605
rect 404262 534692 404268 534744
rect 404320 534732 404326 534744
rect 473906 534732 473912 534744
rect 404320 534704 473912 534732
rect 404320 534692 404326 534704
rect 473906 534692 473912 534704
rect 473964 534692 473970 534744
rect 331490 534664 331496 534676
rect 331451 534636 331496 534664
rect 331490 534624 331496 534636
rect 331548 534624 331554 534676
rect 331306 534460 331312 534472
rect 331219 534432 331312 534460
rect 331306 534420 331312 534432
rect 331364 534460 331370 534472
rect 334894 534460 334900 534472
rect 331364 534432 334900 534460
rect 331364 534420 331370 534432
rect 334894 534420 334900 534432
rect 334952 534420 334958 534472
rect 331490 534284 331496 534336
rect 331548 534324 331554 534336
rect 402974 534324 402980 534336
rect 331548 534296 402980 534324
rect 331548 534284 331554 534296
rect 402974 534284 402980 534296
rect 403032 534324 403038 534336
rect 404262 534324 404268 534336
rect 403032 534296 404268 534324
rect 403032 534284 403038 534296
rect 404262 534284 404268 534296
rect 404320 534284 404326 534336
rect 136177 533987 136235 533993
rect 136177 533953 136189 533987
rect 136223 533984 136235 533987
rect 361482 533984 361488 533996
rect 136223 533956 361488 533984
rect 136223 533953 136235 533956
rect 136177 533947 136235 533953
rect 361482 533944 361488 533956
rect 361540 533944 361546 533996
rect 4522 533740 4528 533792
rect 4580 533780 4586 533792
rect 136085 533783 136143 533789
rect 136085 533780 136097 533783
rect 4580 533752 136097 533780
rect 4580 533740 4586 533752
rect 136085 533749 136097 533752
rect 136131 533780 136143 533783
rect 430758 533780 430764 533792
rect 136131 533752 430764 533780
rect 136131 533749 136143 533752
rect 136085 533743 136143 533749
rect 430758 533740 430764 533752
rect 430816 533740 430822 533792
rect 342438 531604 342444 531616
rect 342399 531576 342444 531604
rect 342438 531564 342444 531576
rect 342496 531564 342502 531616
rect 355594 529020 355600 529032
rect 355507 528992 355600 529020
rect 355594 528980 355600 528992
rect 355652 529020 355658 529032
rect 417970 529020 417976 529032
rect 355652 528992 417976 529020
rect 355652 528980 355658 528992
rect 417970 528980 417976 528992
rect 418028 528980 418034 529032
rect 355502 528884 355508 528896
rect 355463 528856 355508 528884
rect 355502 528844 355508 528856
rect 355560 528844 355566 528896
rect 121822 528504 121828 528556
rect 121880 528544 121886 528556
rect 495434 528544 495440 528556
rect 121880 528516 495440 528544
rect 121880 528504 121886 528516
rect 495434 528504 495440 528516
rect 495492 528504 495498 528556
rect 81342 528300 81348 528352
rect 81400 528340 81406 528352
rect 91373 528343 91431 528349
rect 91373 528340 91385 528343
rect 81400 528312 91385 528340
rect 81400 528300 81406 528312
rect 91373 528309 91385 528312
rect 91419 528309 91431 528343
rect 91373 528303 91431 528309
rect 12986 527932 12992 527944
rect 12947 527904 12992 527932
rect 12986 527892 12992 527904
rect 13044 527892 13050 527944
rect 353938 527932 353944 527944
rect 353899 527904 353944 527932
rect 353938 527892 353944 527904
rect 353996 527892 354002 527944
rect 12710 527864 12716 527876
rect 12768 527873 12774 527876
rect 12680 527836 12716 527864
rect 12710 527824 12716 527836
rect 12768 527827 12780 527873
rect 12768 527824 12774 527827
rect 11609 527799 11667 527805
rect 11609 527765 11621 527799
rect 11655 527796 11667 527799
rect 417786 527796 417792 527808
rect 11655 527768 417792 527796
rect 11655 527765 11667 527768
rect 11609 527759 11667 527765
rect 417786 527756 417792 527768
rect 417844 527756 417850 527808
rect 112530 527416 112536 527468
rect 112588 527456 112594 527468
rect 376766 527459 376824 527465
rect 376766 527456 376778 527459
rect 112588 527428 376778 527456
rect 112588 527416 112594 527428
rect 376766 527425 376778 527428
rect 376812 527425 376824 527459
rect 376766 527419 376824 527425
rect 377033 527459 377091 527465
rect 377033 527425 377045 527459
rect 377079 527456 377091 527459
rect 380618 527456 380624 527468
rect 377079 527428 380624 527456
rect 377079 527425 377091 527428
rect 377033 527419 377091 527425
rect 380618 527416 380624 527428
rect 380676 527416 380682 527468
rect 375650 527252 375656 527264
rect 375611 527224 375656 527252
rect 375650 527212 375656 527224
rect 375708 527212 375714 527264
rect 380618 527144 380624 527196
rect 380676 527184 380682 527196
rect 383654 527184 383660 527196
rect 380676 527156 383660 527184
rect 380676 527144 380682 527156
rect 383654 527144 383660 527156
rect 383712 527144 383718 527196
rect 121089 526371 121147 526377
rect 121089 526337 121101 526371
rect 121135 526368 121147 526371
rect 273622 526368 273628 526380
rect 121135 526340 273628 526368
rect 121135 526337 121147 526340
rect 121089 526331 121147 526337
rect 273622 526328 273628 526340
rect 273680 526328 273686 526380
rect 120994 526164 121000 526176
rect 120955 526136 121000 526164
rect 120994 526124 121000 526136
rect 121052 526164 121058 526176
rect 158714 526164 158720 526176
rect 121052 526136 158720 526164
rect 121052 526124 121058 526136
rect 158714 526124 158720 526136
rect 158772 526124 158778 526176
rect 262766 525280 262772 525292
rect 262727 525252 262772 525280
rect 262766 525240 262772 525252
rect 262824 525240 262830 525292
rect 351472 525252 354674 525280
rect 351472 525224 351500 525252
rect 262490 525212 262496 525224
rect 262451 525184 262496 525212
rect 262490 525172 262496 525184
rect 262548 525172 262554 525224
rect 262674 525212 262680 525224
rect 262635 525184 262680 525212
rect 262674 525172 262680 525184
rect 262732 525172 262738 525224
rect 290826 525212 290832 525224
rect 267706 525184 290832 525212
rect 262508 525144 262536 525172
rect 267706 525144 267734 525184
rect 290826 525172 290832 525184
rect 290884 525172 290890 525224
rect 351454 525212 351460 525224
rect 351415 525184 351460 525212
rect 351454 525172 351460 525184
rect 351512 525172 351518 525224
rect 351730 525212 351736 525224
rect 351691 525184 351736 525212
rect 351730 525172 351736 525184
rect 351788 525172 351794 525224
rect 354646 525212 354674 525252
rect 452102 525212 452108 525224
rect 354646 525184 452108 525212
rect 452102 525172 452108 525184
rect 452160 525172 452166 525224
rect 262508 525116 267734 525144
rect 12345 525079 12403 525085
rect 12345 525045 12357 525079
rect 12391 525076 12403 525079
rect 15286 525076 15292 525088
rect 12391 525048 15292 525076
rect 12391 525045 12403 525048
rect 12345 525039 12403 525045
rect 15286 525036 15292 525048
rect 15344 525076 15350 525088
rect 153470 525076 153476 525088
rect 15344 525048 153476 525076
rect 15344 525036 15350 525048
rect 153470 525036 153476 525048
rect 153528 525036 153534 525088
rect 263137 525079 263195 525085
rect 263137 525045 263149 525079
rect 263183 525076 263195 525079
rect 350905 525079 350963 525085
rect 350905 525076 350917 525079
rect 263183 525048 350917 525076
rect 263183 525045 263195 525048
rect 263137 525039 263195 525045
rect 350905 525045 350917 525048
rect 350951 525045 350963 525079
rect 350905 525039 350963 525045
rect 158622 524804 158628 524816
rect 10888 524776 158628 524804
rect 10888 524745 10916 524776
rect 158622 524764 158628 524776
rect 158680 524764 158686 524816
rect 10873 524739 10931 524745
rect 10873 524705 10885 524739
rect 10919 524705 10931 524739
rect 10873 524699 10931 524705
rect 11517 524739 11575 524745
rect 11517 524705 11529 524739
rect 11563 524736 11575 524739
rect 75914 524736 75920 524748
rect 11563 524708 75920 524736
rect 11563 524705 11575 524708
rect 11517 524699 11575 524705
rect 75914 524696 75920 524708
rect 75972 524696 75978 524748
rect 350905 524739 350963 524745
rect 350905 524705 350917 524739
rect 350951 524736 350963 524739
rect 351549 524739 351607 524745
rect 351549 524736 351561 524739
rect 350951 524708 351561 524736
rect 350951 524705 350963 524708
rect 350905 524699 350963 524705
rect 351549 524705 351561 524708
rect 351595 524705 351607 524739
rect 351730 524736 351736 524748
rect 351691 524708 351736 524736
rect 351549 524699 351607 524705
rect 351730 524696 351736 524708
rect 351788 524696 351794 524748
rect 11241 524671 11299 524677
rect 11241 524637 11253 524671
rect 11287 524637 11299 524671
rect 11241 524631 11299 524637
rect 11701 524671 11759 524677
rect 11701 524637 11713 524671
rect 11747 524668 11759 524671
rect 11747 524640 16574 524668
rect 11747 524637 11759 524640
rect 11701 524631 11759 524637
rect 11256 524600 11284 524631
rect 12345 524603 12403 524609
rect 12345 524600 12357 524603
rect 11256 524572 12357 524600
rect 12345 524569 12357 524572
rect 12391 524569 12403 524603
rect 16546 524600 16574 524640
rect 27430 524600 27436 524612
rect 16546 524572 27436 524600
rect 12345 524563 12403 524569
rect 27430 524560 27436 524572
rect 27488 524560 27494 524612
rect 157518 524560 157524 524612
rect 157576 524600 157582 524612
rect 351457 524603 351515 524609
rect 351457 524600 351469 524603
rect 157576 524572 351469 524600
rect 157576 524560 157582 524572
rect 351457 524569 351469 524572
rect 351503 524569 351515 524603
rect 351457 524563 351515 524569
rect 11422 524532 11428 524544
rect 11383 524504 11428 524532
rect 11422 524492 11428 524504
rect 11480 524492 11486 524544
rect 113082 524492 113088 524544
rect 113140 524532 113146 524544
rect 351089 524535 351147 524541
rect 351089 524532 351101 524535
rect 113140 524504 351101 524532
rect 113140 524492 113146 524504
rect 351089 524501 351101 524504
rect 351135 524501 351147 524535
rect 351089 524495 351147 524501
rect 291102 518752 291108 518764
rect 291063 518724 291108 518752
rect 291102 518712 291108 518724
rect 291160 518712 291166 518764
rect 289814 518644 289820 518696
rect 289872 518684 289878 518696
rect 291197 518687 291255 518693
rect 291197 518684 291209 518687
rect 289872 518656 291209 518684
rect 289872 518644 289878 518656
rect 291197 518653 291209 518656
rect 291243 518653 291255 518687
rect 291197 518647 291255 518653
rect 291289 518687 291347 518693
rect 291289 518653 291301 518687
rect 291335 518653 291347 518687
rect 291289 518647 291347 518653
rect 290826 518576 290832 518628
rect 290884 518616 290890 518628
rect 291304 518616 291332 518647
rect 290884 518588 291332 518616
rect 290884 518576 290890 518588
rect 244918 518508 244924 518560
rect 244976 518548 244982 518560
rect 290737 518551 290795 518557
rect 290737 518548 290749 518551
rect 244976 518520 290749 518548
rect 244976 518508 244982 518520
rect 290737 518517 290749 518520
rect 290783 518517 290795 518551
rect 290737 518511 290795 518517
rect 319898 514876 319904 514888
rect 319859 514848 319904 514876
rect 319898 514836 319904 514848
rect 319956 514876 319962 514888
rect 435082 514876 435088 514888
rect 319956 514848 435088 514876
rect 319956 514836 319962 514848
rect 435082 514836 435088 514848
rect 435140 514836 435146 514888
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 14458 514808 14464 514820
rect 3384 514780 14464 514808
rect 3384 514768 3390 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 319806 514808 319812 514820
rect 319767 514780 319812 514808
rect 319806 514768 319812 514780
rect 319864 514768 319870 514820
rect 92017 514403 92075 514409
rect 92017 514369 92029 514403
rect 92063 514400 92075 514403
rect 309686 514400 309692 514412
rect 92063 514372 309692 514400
rect 92063 514369 92075 514372
rect 92017 514363 92075 514369
rect 309686 514360 309692 514372
rect 309744 514360 309750 514412
rect 405737 514403 405795 514409
rect 405737 514400 405749 514403
rect 393286 514372 405749 514400
rect 267642 514292 267648 514344
rect 267700 514332 267706 514344
rect 393286 514332 393314 514372
rect 405737 514369 405749 514372
rect 405783 514369 405795 514403
rect 405737 514363 405795 514369
rect 405826 514332 405832 514344
rect 267700 514304 393314 514332
rect 405787 514304 405832 514332
rect 267700 514292 267706 514304
rect 405826 514292 405832 514304
rect 405884 514292 405890 514344
rect 406010 514292 406016 514344
rect 406068 514332 406074 514344
rect 409598 514332 409604 514344
rect 406068 514304 409604 514332
rect 406068 514292 406074 514304
rect 409598 514292 409604 514304
rect 409656 514292 409662 514344
rect 92109 514199 92167 514205
rect 92109 514165 92121 514199
rect 92155 514196 92167 514199
rect 157242 514196 157248 514208
rect 92155 514168 157248 514196
rect 92155 514165 92167 514168
rect 92109 514159 92167 514165
rect 157242 514156 157248 514168
rect 157300 514156 157306 514208
rect 405366 514196 405372 514208
rect 405327 514168 405372 514196
rect 405366 514156 405372 514168
rect 405424 514156 405430 514208
rect 46201 513995 46259 514001
rect 46201 513961 46213 513995
rect 46247 513992 46259 513995
rect 328454 513992 328460 514004
rect 46247 513964 328460 513992
rect 46247 513961 46259 513964
rect 46201 513955 46259 513961
rect 328454 513952 328460 513964
rect 328512 513952 328518 514004
rect 26206 513828 55214 513856
rect 24397 513791 24455 513797
rect 24397 513757 24409 513791
rect 24443 513788 24455 513791
rect 26206 513788 26234 513828
rect 45925 513791 45983 513797
rect 45925 513788 45937 513791
rect 24443 513760 26234 513788
rect 45526 513760 45937 513788
rect 24443 513757 24455 513760
rect 24397 513751 24455 513757
rect 7834 513680 7840 513732
rect 7892 513720 7898 513732
rect 45526 513720 45554 513760
rect 45925 513757 45937 513760
rect 45971 513757 45983 513791
rect 45925 513751 45983 513757
rect 46014 513748 46020 513800
rect 46072 513788 46078 513800
rect 55186 513788 55214 513828
rect 260650 513816 260656 513868
rect 260708 513856 260714 513868
rect 276934 513856 276940 513868
rect 260708 513828 276940 513856
rect 260708 513816 260714 513828
rect 276934 513816 276940 513828
rect 276992 513816 276998 513868
rect 410518 513788 410524 513800
rect 46072 513760 46117 513788
rect 55186 513760 260604 513788
rect 46072 513748 46078 513760
rect 46198 513720 46204 513732
rect 7892 513692 45554 513720
rect 46159 513692 46204 513720
rect 7892 513680 7898 513692
rect 46198 513680 46204 513692
rect 46256 513680 46262 513732
rect 177022 513680 177028 513732
rect 177080 513720 177086 513732
rect 260386 513723 260444 513729
rect 260386 513720 260398 513723
rect 177080 513692 260398 513720
rect 177080 513680 177086 513692
rect 260386 513689 260398 513692
rect 260432 513689 260444 513723
rect 260576 513720 260604 513760
rect 267706 513760 410524 513788
rect 267706 513720 267734 513760
rect 410518 513748 410524 513760
rect 410576 513748 410582 513800
rect 260576 513692 267734 513720
rect 260386 513683 260444 513689
rect 45738 513652 45744 513664
rect 45699 513624 45744 513652
rect 45738 513612 45744 513624
rect 45796 513612 45802 513664
rect 259178 513612 259184 513664
rect 259236 513652 259242 513664
rect 259273 513655 259331 513661
rect 259273 513652 259285 513655
rect 259236 513624 259285 513652
rect 259236 513612 259242 513624
rect 259273 513621 259285 513624
rect 259319 513621 259331 513655
rect 259273 513615 259331 513621
rect 317322 510932 317328 510944
rect 317283 510904 317328 510932
rect 317322 510892 317328 510904
rect 317380 510892 317386 510944
rect 8018 509260 8024 509312
rect 8076 509300 8082 509312
rect 495434 509300 495440 509312
rect 8076 509272 495440 509300
rect 8076 509260 8082 509272
rect 495434 509260 495440 509272
rect 495492 509260 495498 509312
rect 326338 508008 326344 508020
rect 326251 507980 326344 508008
rect 326338 507968 326344 507980
rect 326396 507968 326402 508020
rect 326356 507940 326384 507968
rect 496354 507940 496360 507952
rect 326356 507912 496360 507940
rect 496354 507900 496360 507912
rect 496412 507900 496418 507952
rect 59170 507832 59176 507884
rect 59228 507872 59234 507884
rect 325217 507875 325275 507881
rect 325217 507872 325229 507875
rect 59228 507844 325229 507872
rect 59228 507832 59234 507844
rect 325217 507841 325229 507844
rect 325263 507841 325275 507875
rect 426618 507872 426624 507884
rect 426579 507844 426624 507872
rect 325217 507835 325275 507841
rect 426618 507832 426624 507844
rect 426676 507832 426682 507884
rect 426802 507872 426808 507884
rect 426763 507844 426808 507872
rect 426802 507832 426808 507844
rect 426860 507832 426866 507884
rect 324958 507804 324964 507816
rect 324919 507776 324964 507804
rect 324958 507764 324964 507776
rect 325016 507764 325022 507816
rect 326264 507708 335354 507736
rect 324958 507628 324964 507680
rect 325016 507668 325022 507680
rect 326264 507668 326292 507708
rect 325016 507640 326292 507668
rect 335326 507668 335354 507708
rect 383930 507668 383936 507680
rect 335326 507640 383936 507668
rect 325016 507628 325022 507640
rect 383930 507628 383936 507640
rect 383988 507628 383994 507680
rect 426894 507668 426900 507680
rect 426855 507640 426900 507668
rect 426894 507628 426900 507640
rect 426952 507628 426958 507680
rect 247678 507464 247684 507476
rect 247639 507436 247684 507464
rect 247678 507424 247684 507436
rect 247736 507424 247742 507476
rect 248509 507399 248567 507405
rect 248509 507396 248521 507399
rect 247880 507368 248521 507396
rect 247586 507260 247592 507272
rect 247547 507232 247592 507260
rect 247586 507220 247592 507232
rect 247644 507220 247650 507272
rect 247880 507269 247908 507368
rect 248509 507365 248521 507368
rect 248555 507365 248567 507399
rect 248509 507359 248567 507365
rect 248386 507300 258074 507328
rect 247865 507263 247923 507269
rect 247865 507229 247877 507263
rect 247911 507229 247923 507263
rect 247865 507223 247923 507229
rect 247957 507263 248015 507269
rect 247957 507229 247969 507263
rect 248003 507260 248015 507263
rect 248386 507260 248414 507300
rect 248003 507232 248414 507260
rect 250073 507263 250131 507269
rect 248003 507229 248015 507232
rect 247957 507223 248015 507229
rect 250073 507229 250085 507263
rect 250119 507229 250131 507263
rect 258046 507260 258074 507300
rect 496354 507260 496360 507272
rect 258046 507232 496360 507260
rect 250073 507223 250131 507229
rect 41782 507152 41788 507204
rect 41840 507192 41846 507204
rect 248877 507195 248935 507201
rect 248877 507192 248889 507195
rect 41840 507164 248889 507192
rect 41840 507152 41846 507164
rect 248877 507161 248889 507164
rect 248923 507161 248935 507195
rect 250088 507192 250116 507223
rect 496354 507220 496360 507232
rect 496412 507220 496418 507272
rect 250257 507195 250315 507201
rect 250257 507192 250269 507195
rect 250088 507164 250269 507192
rect 248877 507155 248935 507161
rect 250257 507161 250269 507164
rect 250303 507192 250315 507195
rect 373810 507192 373816 507204
rect 250303 507164 373816 507192
rect 250303 507161 250315 507164
rect 250257 507155 250315 507161
rect 373810 507152 373816 507164
rect 373868 507152 373874 507204
rect 248138 507124 248144 507136
rect 248099 507096 248144 507124
rect 248138 507084 248144 507096
rect 248196 507084 248202 507136
rect 248509 506923 248567 506929
rect 248509 506889 248521 506923
rect 248555 506920 248567 506923
rect 248785 506923 248843 506929
rect 248785 506920 248797 506923
rect 248555 506892 248797 506920
rect 248555 506889 248567 506892
rect 248509 506883 248567 506889
rect 248785 506889 248797 506892
rect 248831 506889 248843 506923
rect 248785 506883 248843 506889
rect 249245 506787 249303 506793
rect 249245 506753 249257 506787
rect 249291 506784 249303 506787
rect 250257 506787 250315 506793
rect 250257 506784 250269 506787
rect 249291 506756 250269 506784
rect 249291 506753 249303 506756
rect 249245 506747 249303 506753
rect 250257 506753 250269 506756
rect 250303 506753 250315 506787
rect 250257 506747 250315 506753
rect 3142 505112 3148 505164
rect 3200 505152 3206 505164
rect 349798 505152 349804 505164
rect 3200 505124 349804 505152
rect 3200 505112 3206 505124
rect 349798 505112 349804 505124
rect 349856 505112 349862 505164
rect 383933 504611 383991 504617
rect 383933 504577 383945 504611
rect 383979 504608 383991 504611
rect 384022 504608 384028 504620
rect 383979 504580 384028 504608
rect 383979 504577 383991 504580
rect 383933 504571 383991 504577
rect 384022 504568 384028 504580
rect 384080 504608 384086 504620
rect 406562 504608 406568 504620
rect 384080 504580 406568 504608
rect 384080 504568 384086 504580
rect 406562 504568 406568 504580
rect 406620 504568 406626 504620
rect 383838 504404 383844 504416
rect 383751 504376 383844 504404
rect 383838 504364 383844 504376
rect 383896 504404 383902 504416
rect 443086 504404 443092 504416
rect 383896 504376 443092 504404
rect 383896 504364 383902 504376
rect 443086 504364 443092 504376
rect 443144 504364 443150 504416
rect 406562 503684 406568 503736
rect 406620 503724 406626 503736
rect 464154 503724 464160 503736
rect 406620 503696 464160 503724
rect 406620 503684 406626 503696
rect 464154 503684 464160 503696
rect 464212 503684 464218 503736
rect 116765 502231 116823 502237
rect 116765 502197 116777 502231
rect 116811 502228 116823 502231
rect 153838 502228 153844 502240
rect 116811 502200 153844 502228
rect 116811 502197 116823 502200
rect 116765 502191 116823 502197
rect 153838 502188 153844 502200
rect 153896 502188 153902 502240
rect 421006 500828 421012 500880
rect 421064 500828 421070 500880
rect 420730 500800 420736 500812
rect 420691 500772 420736 500800
rect 420730 500760 420736 500772
rect 420788 500760 420794 500812
rect 420914 500732 420920 500744
rect 420875 500704 420920 500732
rect 420914 500692 420920 500704
rect 420972 500692 420978 500744
rect 421024 500741 421052 500828
rect 421009 500735 421067 500741
rect 421009 500701 421021 500735
rect 421055 500701 421067 500735
rect 421009 500695 421067 500701
rect 421116 500704 422294 500732
rect 420546 500664 420552 500676
rect 420507 500636 420552 500664
rect 420546 500624 420552 500636
rect 420604 500624 420610 500676
rect 420638 500624 420644 500676
rect 420696 500664 420702 500676
rect 421116 500664 421144 500704
rect 420696 500636 421144 500664
rect 421193 500667 421251 500673
rect 420696 500624 420702 500636
rect 421193 500633 421205 500667
rect 421239 500633 421251 500667
rect 422266 500664 422294 500704
rect 481818 500664 481824 500676
rect 422266 500636 481824 500664
rect 421193 500627 421251 500633
rect 369118 500556 369124 500608
rect 369176 500596 369182 500608
rect 421208 500596 421236 500627
rect 481818 500624 481824 500636
rect 481876 500624 481882 500676
rect 369176 500568 421236 500596
rect 369176 500556 369182 500568
rect 190362 500052 190368 500064
rect 190323 500024 190368 500052
rect 190362 500012 190368 500024
rect 190420 500012 190426 500064
rect 208213 498151 208271 498157
rect 208213 498117 208225 498151
rect 208259 498148 208271 498151
rect 208302 498148 208308 498160
rect 208259 498120 208308 498148
rect 208259 498117 208271 498120
rect 208213 498111 208271 498117
rect 208302 498108 208308 498120
rect 208360 498108 208366 498160
rect 208397 498151 208455 498157
rect 208397 498117 208409 498151
rect 208443 498148 208455 498151
rect 208443 498120 209774 498148
rect 208443 498117 208455 498120
rect 208397 498111 208455 498117
rect 208578 498080 208584 498092
rect 208539 498052 208584 498080
rect 208578 498040 208584 498052
rect 208636 498040 208642 498092
rect 209746 498080 209774 498120
rect 233786 498080 233792 498092
rect 209746 498052 233792 498080
rect 233786 498040 233792 498052
rect 233844 498040 233850 498092
rect 208302 497836 208308 497888
rect 208360 497876 208366 497888
rect 331582 497876 331588 497888
rect 208360 497848 331588 497876
rect 208360 497836 208366 497848
rect 331582 497836 331588 497848
rect 331640 497836 331646 497888
rect 2774 496952 2780 497004
rect 2832 496992 2838 497004
rect 5350 496992 5356 497004
rect 2832 496964 5356 496992
rect 2832 496952 2838 496964
rect 5350 496952 5356 496964
rect 5408 496952 5414 497004
rect 256789 496451 256847 496457
rect 256789 496448 256801 496451
rect 255608 496420 256801 496448
rect 255608 496392 255636 496420
rect 256789 496417 256801 496420
rect 256835 496417 256847 496451
rect 256789 496411 256847 496417
rect 255590 496380 255596 496392
rect 255551 496352 255596 496380
rect 255590 496340 255596 496352
rect 255648 496340 255654 496392
rect 256053 496383 256111 496389
rect 256053 496349 256065 496383
rect 256099 496380 256111 496383
rect 256329 496383 256387 496389
rect 256329 496380 256341 496383
rect 256099 496352 256341 496380
rect 256099 496349 256111 496352
rect 256053 496343 256111 496349
rect 256329 496349 256341 496352
rect 256375 496349 256387 496383
rect 256329 496343 256387 496349
rect 255777 496247 255835 496253
rect 255777 496213 255789 496247
rect 255823 496244 255835 496247
rect 351454 496244 351460 496256
rect 255823 496216 351460 496244
rect 255823 496213 255835 496216
rect 255777 496207 255835 496213
rect 351454 496204 351460 496216
rect 351512 496204 351518 496256
rect 423582 496108 423588 496120
rect 383626 496080 423588 496108
rect 255869 496043 255927 496049
rect 255869 496009 255881 496043
rect 255915 496040 255927 496043
rect 256053 496043 256111 496049
rect 256053 496040 256065 496043
rect 255915 496012 256065 496040
rect 255915 496009 255927 496012
rect 255869 496003 255927 496009
rect 256053 496009 256065 496012
rect 256099 496009 256111 496043
rect 256053 496003 256111 496009
rect 255700 495944 258074 495972
rect 255700 495916 255728 495944
rect 255682 495904 255688 495916
rect 255643 495876 255688 495904
rect 255682 495864 255688 495876
rect 255740 495864 255746 495916
rect 256329 495907 256387 495913
rect 256329 495873 256341 495907
rect 256375 495873 256387 495907
rect 258046 495904 258074 495944
rect 380710 495904 380716 495916
rect 258046 495876 380716 495904
rect 256329 495867 256387 495873
rect 255590 495796 255596 495848
rect 255648 495836 255654 495848
rect 256344 495836 256372 495867
rect 380710 495864 380716 495876
rect 380768 495904 380774 495916
rect 383626 495904 383654 496080
rect 423582 496068 423588 496080
rect 423640 496068 423646 496120
rect 380768 495876 383654 495904
rect 380768 495864 380774 495876
rect 255648 495808 256372 495836
rect 257157 495839 257215 495845
rect 255648 495796 255654 495808
rect 257157 495805 257169 495839
rect 257203 495836 257215 495839
rect 290274 495836 290280 495848
rect 257203 495808 290280 495836
rect 257203 495805 257215 495808
rect 257157 495799 257215 495805
rect 290274 495796 290280 495808
rect 290332 495796 290338 495848
rect 6454 494572 6460 494624
rect 6512 494612 6518 494624
rect 204901 494615 204959 494621
rect 204901 494612 204913 494615
rect 6512 494584 204913 494612
rect 6512 494572 6518 494584
rect 204901 494581 204913 494584
rect 204947 494581 204959 494615
rect 204901 494575 204959 494581
rect 3694 494164 3700 494216
rect 3752 494204 3758 494216
rect 229097 494207 229155 494213
rect 229097 494204 229109 494207
rect 3752 494176 229109 494204
rect 3752 494164 3758 494176
rect 229097 494173 229109 494176
rect 229143 494173 229155 494207
rect 229097 494167 229155 494173
rect 29638 493144 29644 493196
rect 29696 493184 29702 493196
rect 32125 493187 32183 493193
rect 32125 493184 32137 493187
rect 29696 493156 32137 493184
rect 29696 493144 29702 493156
rect 32125 493153 32137 493156
rect 32171 493184 32183 493187
rect 93762 493184 93768 493196
rect 32171 493156 93768 493184
rect 32171 493153 32183 493156
rect 32125 493147 32183 493153
rect 93762 493144 93768 493156
rect 93820 493144 93826 493196
rect 32306 493048 32312 493060
rect 32267 493020 32312 493048
rect 32306 493008 32312 493020
rect 32364 493008 32370 493060
rect 32398 492940 32404 492992
rect 32456 492980 32462 492992
rect 32766 492980 32772 492992
rect 32456 492952 32501 492980
rect 32727 492952 32772 492980
rect 32456 492940 32462 492952
rect 32766 492940 32772 492952
rect 32824 492940 32830 492992
rect 276934 492192 276940 492244
rect 276992 492232 276998 492244
rect 276992 492204 287054 492232
rect 276992 492192 276998 492204
rect 278317 492167 278375 492173
rect 278317 492133 278329 492167
rect 278363 492164 278375 492167
rect 278685 492167 278743 492173
rect 278685 492164 278697 492167
rect 278363 492136 278697 492164
rect 278363 492133 278375 492136
rect 278317 492127 278375 492133
rect 278685 492133 278697 492136
rect 278731 492133 278743 492167
rect 278685 492127 278743 492133
rect 276934 492096 276940 492108
rect 276895 492068 276940 492096
rect 276934 492056 276940 492068
rect 276992 492056 276998 492108
rect 208486 492028 208492 492040
rect 208447 492000 208492 492028
rect 208486 491988 208492 492000
rect 208544 492028 208550 492040
rect 237374 492028 237380 492040
rect 208544 492000 237380 492028
rect 208544 491988 208550 492000
rect 237374 491988 237380 492000
rect 237432 491988 237438 492040
rect 287026 492028 287054 492204
rect 324958 492028 324964 492040
rect 277044 492000 278728 492028
rect 287026 492000 324964 492028
rect 208244 491963 208302 491969
rect 208244 491929 208256 491963
rect 208290 491960 208302 491963
rect 277044 491960 277072 492000
rect 208290 491932 277072 491960
rect 277204 491963 277262 491969
rect 208290 491929 208302 491932
rect 208244 491923 208302 491929
rect 277204 491929 277216 491963
rect 277250 491960 277262 491963
rect 277302 491960 277308 491972
rect 277250 491932 277308 491960
rect 277250 491929 277262 491932
rect 277204 491923 277262 491929
rect 277302 491920 277308 491932
rect 277360 491920 277366 491972
rect 278700 491960 278728 492000
rect 324958 491988 324964 492000
rect 325016 491988 325022 492040
rect 384298 491960 384304 491972
rect 278240 491932 278544 491960
rect 278700 491932 384304 491960
rect 207106 491892 207112 491904
rect 207067 491864 207112 491892
rect 207106 491852 207112 491864
rect 207164 491892 207170 491904
rect 278240 491892 278268 491932
rect 207164 491864 278268 491892
rect 278516 491892 278544 491932
rect 384298 491920 384304 491932
rect 384356 491920 384362 491972
rect 429286 491892 429292 491904
rect 278516 491864 429292 491892
rect 207164 491852 207170 491864
rect 429286 491852 429292 491864
rect 429344 491852 429350 491904
rect 277302 491648 277308 491700
rect 277360 491688 277366 491700
rect 378778 491688 378784 491700
rect 277360 491660 378784 491688
rect 277360 491648 277366 491660
rect 378778 491648 378784 491660
rect 378836 491648 378842 491700
rect 278685 491623 278743 491629
rect 278685 491589 278697 491623
rect 278731 491620 278743 491623
rect 367002 491620 367008 491632
rect 278731 491592 367008 491620
rect 278731 491589 278743 491592
rect 278685 491583 278743 491589
rect 367002 491580 367008 491592
rect 367060 491580 367066 491632
rect 237374 489812 237380 489864
rect 237432 489852 237438 489864
rect 238202 489852 238208 489864
rect 237432 489824 238208 489852
rect 237432 489812 237438 489824
rect 238202 489812 238208 489824
rect 238260 489852 238266 489864
rect 248049 489855 248107 489861
rect 248049 489852 248061 489855
rect 238260 489824 248061 489852
rect 238260 489812 238266 489824
rect 248049 489821 248061 489824
rect 248095 489852 248107 489855
rect 276934 489852 276940 489864
rect 248095 489824 276940 489852
rect 248095 489821 248107 489824
rect 248049 489815 248107 489821
rect 276934 489812 276940 489824
rect 276992 489812 276998 489864
rect 412910 489852 412916 489864
rect 412823 489824 412916 489852
rect 412910 489812 412916 489824
rect 412968 489852 412974 489864
rect 432506 489852 432512 489864
rect 412968 489824 432512 489852
rect 412968 489812 412974 489824
rect 432506 489812 432512 489824
rect 432564 489812 432570 489864
rect 248322 489793 248328 489796
rect 248316 489784 248328 489793
rect 248283 489756 248328 489784
rect 248316 489747 248328 489756
rect 248322 489744 248328 489747
rect 248380 489744 248386 489796
rect 413158 489787 413216 489793
rect 413158 489784 413170 489787
rect 393286 489756 413170 489784
rect 249426 489716 249432 489728
rect 249387 489688 249432 489716
rect 249426 489676 249432 489688
rect 249484 489676 249490 489728
rect 27522 489472 27528 489524
rect 27580 489512 27586 489524
rect 393286 489512 393314 489756
rect 413158 489753 413170 489756
rect 413204 489753 413216 489787
rect 413158 489747 413216 489753
rect 414290 489716 414296 489728
rect 414251 489688 414296 489716
rect 414290 489676 414296 489688
rect 414348 489716 414354 489728
rect 423950 489716 423956 489728
rect 414348 489688 423956 489716
rect 414348 489676 414354 489688
rect 423950 489676 423956 489688
rect 424008 489676 424014 489728
rect 27580 489484 393314 489512
rect 27580 489472 27586 489484
rect 470042 489172 470048 489184
rect 470003 489144 470048 489172
rect 470042 489132 470048 489144
rect 470100 489132 470106 489184
rect 21453 487339 21511 487345
rect 21453 487305 21465 487339
rect 21499 487336 21511 487339
rect 21634 487336 21640 487348
rect 21499 487308 21640 487336
rect 21499 487305 21511 487308
rect 21453 487299 21511 487305
rect 21634 487296 21640 487308
rect 21692 487296 21698 487348
rect 9582 487228 9588 487280
rect 9640 487268 9646 487280
rect 20993 487271 21051 487277
rect 20993 487268 21005 487271
rect 9640 487240 21005 487268
rect 9640 487228 9646 487240
rect 20993 487237 21005 487240
rect 21039 487237 21051 487271
rect 20993 487231 21051 487237
rect 237650 487228 237656 487280
rect 237708 487268 237714 487280
rect 417513 487271 417571 487277
rect 417513 487268 417525 487271
rect 237708 487240 417525 487268
rect 237708 487228 237714 487240
rect 417513 487237 417525 487240
rect 417559 487237 417571 487271
rect 417513 487231 417571 487237
rect 417786 487228 417792 487280
rect 417844 487228 417850 487280
rect 417878 487228 417884 487280
rect 417936 487228 417942 487280
rect 417788 487225 417846 487228
rect 7098 487160 7104 487212
rect 7156 487200 7162 487212
rect 21085 487203 21143 487209
rect 21085 487200 21097 487203
rect 7156 487172 21097 487200
rect 7156 487160 7162 487172
rect 21085 487169 21097 487172
rect 21131 487169 21143 487203
rect 417788 487191 417800 487225
rect 417834 487191 417846 487225
rect 417788 487185 417846 487191
rect 417880 487225 417938 487228
rect 417880 487191 417892 487225
rect 417926 487191 417938 487225
rect 417880 487185 417938 487191
rect 21085 487163 21143 487169
rect 417970 487160 417976 487212
rect 418028 487200 418034 487212
rect 418157 487203 418215 487209
rect 418028 487172 418073 487200
rect 418028 487160 418034 487172
rect 418157 487169 418169 487203
rect 418203 487200 418215 487203
rect 422018 487200 422024 487212
rect 418203 487172 422024 487200
rect 418203 487169 418215 487172
rect 418157 487163 418215 487169
rect 422018 487160 422024 487172
rect 422076 487160 422082 487212
rect 20901 487135 20959 487141
rect 20901 487101 20913 487135
rect 20947 487101 20959 487135
rect 20901 487095 20959 487101
rect 20916 487064 20944 487095
rect 29638 487064 29644 487076
rect 20916 487036 29644 487064
rect 29638 487024 29644 487036
rect 29696 487024 29702 487076
rect 264054 485636 264060 485648
rect 264015 485608 264060 485636
rect 264054 485596 264060 485608
rect 264112 485596 264118 485648
rect 263686 485528 263692 485580
rect 263744 485568 263750 485580
rect 420730 485568 420736 485580
rect 263744 485540 420736 485568
rect 263744 485528 263750 485540
rect 420730 485528 420736 485540
rect 420788 485528 420794 485580
rect 263870 485500 263876 485512
rect 263831 485472 263876 485500
rect 263870 485460 263876 485472
rect 263928 485500 263934 485512
rect 420546 485500 420552 485512
rect 263928 485472 420552 485500
rect 263928 485460 263934 485472
rect 420546 485460 420552 485472
rect 420604 485460 420610 485512
rect 263520 485404 264008 485432
rect 263520 485376 263548 485404
rect 263502 485364 263508 485376
rect 263463 485336 263508 485364
rect 263502 485324 263508 485336
rect 263560 485324 263566 485376
rect 263686 485364 263692 485376
rect 263647 485336 263692 485364
rect 263686 485324 263692 485336
rect 263744 485324 263750 485376
rect 263778 485324 263784 485376
rect 263836 485364 263842 485376
rect 263980 485364 264008 485404
rect 264146 485392 264152 485444
rect 264204 485432 264210 485444
rect 477770 485432 477776 485444
rect 264204 485404 477776 485432
rect 264204 485392 264210 485404
rect 477770 485392 477776 485404
rect 477828 485392 477834 485444
rect 421006 485364 421012 485376
rect 263836 485336 263881 485364
rect 263980 485336 421012 485364
rect 263836 485324 263842 485336
rect 421006 485324 421012 485336
rect 421064 485324 421070 485376
rect 464154 484072 464160 484084
rect 464115 484044 464160 484072
rect 464154 484032 464160 484044
rect 464212 484032 464218 484084
rect 464246 484032 464252 484084
rect 464304 484072 464310 484084
rect 464304 484044 464349 484072
rect 464304 484032 464310 484044
rect 463970 483936 463976 483948
rect 463931 483908 463976 483936
rect 463970 483896 463976 483908
rect 464028 483896 464034 483948
rect 464338 483936 464344 483948
rect 464299 483908 464344 483936
rect 464338 483896 464344 483908
rect 464396 483896 464402 483948
rect 167270 483760 167276 483812
rect 167328 483800 167334 483812
rect 464525 483803 464583 483809
rect 464525 483800 464537 483803
rect 167328 483772 464537 483800
rect 167328 483760 167334 483772
rect 464525 483769 464537 483772
rect 464571 483769 464583 483803
rect 464525 483763 464583 483769
rect 382550 482440 382556 482452
rect 382511 482412 382556 482440
rect 382550 482400 382556 482412
rect 382608 482400 382614 482452
rect 383930 482304 383936 482316
rect 383891 482276 383936 482304
rect 383930 482264 383936 482276
rect 383988 482304 383994 482316
rect 383988 482276 393314 482304
rect 383988 482264 383994 482276
rect 393286 482236 393314 482276
rect 412910 482236 412916 482248
rect 393286 482208 412916 482236
rect 412910 482196 412916 482208
rect 412968 482196 412974 482248
rect 383666 482171 383724 482177
rect 383666 482137 383678 482171
rect 383712 482137 383724 482171
rect 383666 482131 383724 482137
rect 383672 482100 383700 482131
rect 383746 482100 383752 482112
rect 383672 482072 383752 482100
rect 383746 482060 383752 482072
rect 383804 482060 383810 482112
rect 16393 480675 16451 480681
rect 16393 480641 16405 480675
rect 16439 480672 16451 480675
rect 22830 480672 22836 480684
rect 16439 480644 22836 480672
rect 16439 480641 16451 480644
rect 16393 480635 16451 480641
rect 22830 480632 22836 480644
rect 22888 480632 22894 480684
rect 16577 480607 16635 480613
rect 16577 480573 16589 480607
rect 16623 480604 16635 480607
rect 327718 480604 327724 480616
rect 16623 480576 327724 480604
rect 16623 480573 16635 480576
rect 16577 480567 16635 480573
rect 327718 480564 327724 480576
rect 327776 480564 327782 480616
rect 16206 480468 16212 480480
rect 16167 480440 16212 480468
rect 16206 480428 16212 480440
rect 16264 480428 16270 480480
rect 238202 480128 238208 480140
rect 238163 480100 238208 480128
rect 238202 480088 238208 480100
rect 238260 480088 238266 480140
rect 238478 480001 238484 480004
rect 238472 479955 238484 480001
rect 238536 479992 238542 480004
rect 238536 479964 238572 479992
rect 238478 479952 238484 479955
rect 238536 479952 238542 479964
rect 239585 479927 239643 479933
rect 239585 479893 239597 479927
rect 239631 479924 239643 479927
rect 259362 479924 259368 479936
rect 239631 479896 259368 479924
rect 239631 479893 239643 479896
rect 239585 479887 239643 479893
rect 259362 479884 259368 479896
rect 259420 479884 259426 479936
rect 2774 479000 2780 479052
rect 2832 479040 2838 479052
rect 5258 479040 5264 479052
rect 2832 479012 5264 479040
rect 2832 479000 2838 479012
rect 5258 479000 5264 479012
rect 5316 479000 5322 479052
rect 259362 478864 259368 478916
rect 259420 478904 259426 478916
rect 331674 478904 331680 478916
rect 259420 478876 331680 478904
rect 259420 478864 259426 478876
rect 331674 478864 331680 478876
rect 331732 478864 331738 478916
rect 360562 475736 360568 475788
rect 360620 475776 360626 475788
rect 495345 475779 495403 475785
rect 495345 475776 495357 475779
rect 360620 475748 495357 475776
rect 360620 475736 360626 475748
rect 495345 475745 495357 475748
rect 495391 475745 495403 475779
rect 495345 475739 495403 475745
rect 297634 475668 297640 475720
rect 297692 475708 297698 475720
rect 495253 475711 495311 475717
rect 495253 475708 495265 475711
rect 297692 475680 495265 475708
rect 297692 475668 297698 475680
rect 495253 475677 495265 475680
rect 495299 475677 495311 475711
rect 495526 475708 495532 475720
rect 495487 475680 495532 475708
rect 495253 475671 495311 475677
rect 495526 475668 495532 475680
rect 495584 475668 495590 475720
rect 495618 475668 495624 475720
rect 495676 475708 495682 475720
rect 495676 475680 495721 475708
rect 495676 475668 495682 475680
rect 5902 475532 5908 475584
rect 5960 475572 5966 475584
rect 495805 475575 495863 475581
rect 495805 475572 495817 475575
rect 5960 475544 495817 475572
rect 5960 475532 5966 475544
rect 495805 475541 495817 475544
rect 495851 475541 495863 475575
rect 495805 475535 495863 475541
rect 9766 475328 9772 475380
rect 9824 475368 9830 475380
rect 194594 475368 194600 475380
rect 9824 475340 194600 475368
rect 9824 475328 9830 475340
rect 194594 475328 194600 475340
rect 194652 475328 194658 475380
rect 93762 473628 93768 473680
rect 93820 473628 93826 473680
rect 93780 473600 93808 473628
rect 94041 473603 94099 473609
rect 94041 473600 94053 473603
rect 93780 473572 94053 473600
rect 94041 473569 94053 473572
rect 94087 473600 94099 473603
rect 112438 473600 112444 473612
rect 94087 473572 112444 473600
rect 94087 473569 94099 473572
rect 94041 473563 94099 473569
rect 112438 473560 112444 473572
rect 112496 473560 112502 473612
rect 93762 473492 93768 473544
rect 93820 473532 93826 473544
rect 93857 473535 93915 473541
rect 93857 473532 93869 473535
rect 93820 473504 93869 473532
rect 93820 473492 93826 473504
rect 93857 473501 93869 473504
rect 93903 473501 93915 473535
rect 93857 473495 93915 473501
rect 97074 473492 97080 473544
rect 97132 473532 97138 473544
rect 202693 473535 202751 473541
rect 202693 473532 202705 473535
rect 97132 473504 202705 473532
rect 97132 473492 97138 473504
rect 202693 473501 202705 473504
rect 202739 473501 202751 473535
rect 202693 473495 202751 473501
rect 202877 473535 202935 473541
rect 202877 473501 202889 473535
rect 202923 473532 202935 473535
rect 228910 473532 228916 473544
rect 202923 473504 228916 473532
rect 202923 473501 202935 473504
rect 202877 473495 202935 473501
rect 228910 473492 228916 473504
rect 228968 473492 228974 473544
rect 93302 473356 93308 473408
rect 93360 473396 93366 473408
rect 93397 473399 93455 473405
rect 93397 473396 93409 473399
rect 93360 473368 93409 473396
rect 93360 473356 93366 473368
rect 93397 473365 93409 473368
rect 93443 473365 93455 473399
rect 93397 473359 93455 473365
rect 93670 473356 93676 473408
rect 93728 473396 93734 473408
rect 93765 473399 93823 473405
rect 93765 473396 93777 473399
rect 93728 473368 93777 473396
rect 93728 473356 93734 473368
rect 93765 473365 93777 473368
rect 93811 473365 93823 473399
rect 203058 473396 203064 473408
rect 203019 473368 203064 473396
rect 93765 473359 93823 473365
rect 203058 473356 203064 473368
rect 203116 473356 203122 473408
rect 198645 471359 198703 471365
rect 198645 471325 198657 471359
rect 198691 471356 198703 471359
rect 263502 471356 263508 471368
rect 198691 471328 263508 471356
rect 198691 471325 198703 471328
rect 198645 471319 198703 471325
rect 263502 471316 263508 471328
rect 263560 471316 263566 471368
rect 198274 471288 198280 471300
rect 198235 471260 198280 471288
rect 198274 471248 198280 471260
rect 198332 471248 198338 471300
rect 198458 471248 198464 471300
rect 198516 471288 198522 471300
rect 268838 471288 268844 471300
rect 198516 471260 268844 471288
rect 198516 471248 198522 471260
rect 268838 471248 268844 471260
rect 268896 471248 268902 471300
rect 194778 470948 194784 470960
rect 149348 470920 194784 470948
rect 149348 470889 149376 470920
rect 194778 470908 194784 470920
rect 194836 470908 194842 470960
rect 149333 470883 149391 470889
rect 149333 470849 149345 470883
rect 149379 470849 149391 470883
rect 149333 470843 149391 470849
rect 149600 470883 149658 470889
rect 149600 470849 149612 470883
rect 149646 470880 149658 470883
rect 344278 470880 344284 470892
rect 149646 470852 344284 470880
rect 149646 470849 149658 470852
rect 149600 470843 149658 470849
rect 344278 470840 344284 470852
rect 344336 470840 344342 470892
rect 150713 470679 150771 470685
rect 150713 470645 150725 470679
rect 150759 470676 150771 470679
rect 384022 470676 384028 470688
rect 150759 470648 384028 470676
rect 150759 470645 150771 470648
rect 150713 470639 150771 470645
rect 384022 470636 384028 470648
rect 384080 470636 384086 470688
rect 432417 469863 432475 469869
rect 432417 469829 432429 469863
rect 432463 469860 432475 469863
rect 432506 469860 432512 469872
rect 432463 469832 432512 469860
rect 432463 469829 432475 469832
rect 432417 469823 432475 469829
rect 432506 469820 432512 469832
rect 432564 469860 432570 469872
rect 443914 469860 443920 469872
rect 432564 469832 443920 469860
rect 432564 469820 432570 469832
rect 443914 469820 443920 469832
rect 443972 469860 443978 469872
rect 494330 469860 494336 469872
rect 443972 469832 494336 469860
rect 443972 469820 443978 469832
rect 494330 469820 494336 469832
rect 494388 469820 494394 469872
rect 167914 469752 167920 469804
rect 167972 469792 167978 469804
rect 432765 469795 432823 469801
rect 432765 469792 432777 469795
rect 167972 469764 432777 469792
rect 167972 469752 167978 469764
rect 432765 469761 432777 469764
rect 432811 469761 432823 469795
rect 432765 469755 432823 469761
rect 432417 469727 432475 469733
rect 432417 469693 432429 469727
rect 432463 469724 432475 469727
rect 432509 469727 432567 469733
rect 432509 469724 432521 469727
rect 432463 469696 432521 469724
rect 432463 469693 432475 469696
rect 432417 469687 432475 469693
rect 432509 469693 432521 469696
rect 432555 469693 432567 469727
rect 432509 469687 432567 469693
rect 8938 469548 8944 469600
rect 8996 469588 9002 469600
rect 433889 469591 433947 469597
rect 433889 469588 433901 469591
rect 8996 469560 433901 469588
rect 8996 469548 9002 469560
rect 433889 469557 433901 469560
rect 433935 469588 433947 469591
rect 463970 469588 463976 469600
rect 433935 469560 463976 469588
rect 433935 469557 433947 469560
rect 433889 469551 433947 469557
rect 463970 469548 463976 469560
rect 464028 469548 464034 469600
rect 315758 469208 315764 469260
rect 315816 469248 315822 469260
rect 495434 469248 495440 469260
rect 315816 469220 495440 469248
rect 315816 469208 315822 469220
rect 495434 469208 495440 469220
rect 495492 469208 495498 469260
rect 112625 467483 112683 467489
rect 112625 467449 112637 467483
rect 112671 467480 112683 467483
rect 334618 467480 334624 467492
rect 112671 467452 334624 467480
rect 112671 467449 112683 467452
rect 112625 467443 112683 467449
rect 334618 467440 334624 467452
rect 334676 467440 334682 467492
rect 112990 467372 112996 467424
rect 113048 467412 113054 467424
rect 247586 467412 247592 467424
rect 113048 467384 247592 467412
rect 113048 467372 113054 467384
rect 247586 467372 247592 467384
rect 247644 467372 247650 467424
rect 111886 467208 111892 467220
rect 111847 467180 111892 467208
rect 111886 467168 111892 467180
rect 111944 467168 111950 467220
rect 194778 467208 194784 467220
rect 194691 467180 194784 467208
rect 194778 467168 194784 467180
rect 194836 467208 194842 467220
rect 208486 467208 208492 467220
rect 194836 467180 208492 467208
rect 194836 467168 194842 467180
rect 208486 467168 208492 467180
rect 208544 467168 208550 467220
rect 112625 467143 112683 467149
rect 112625 467140 112637 467143
rect 112088 467112 112637 467140
rect 112088 467013 112116 467112
rect 112625 467109 112637 467112
rect 112671 467109 112683 467143
rect 112625 467103 112683 467109
rect 112349 467075 112407 467081
rect 112349 467041 112361 467075
rect 112395 467072 112407 467075
rect 112990 467072 112996 467084
rect 112395 467044 112996 467072
rect 112395 467041 112407 467044
rect 112349 467035 112407 467041
rect 112990 467032 112996 467044
rect 113048 467032 113054 467084
rect 194796 467081 194824 467168
rect 194781 467075 194839 467081
rect 194781 467041 194793 467075
rect 194827 467041 194839 467075
rect 194781 467035 194839 467041
rect 112073 467007 112131 467013
rect 112073 466973 112085 467007
rect 112119 466973 112131 467007
rect 112073 466967 112131 466973
rect 112165 467007 112223 467013
rect 112165 466973 112177 467007
rect 112211 466973 112223 467007
rect 112165 466967 112223 466973
rect 112441 467007 112499 467013
rect 112441 466973 112453 467007
rect 112487 467004 112499 467007
rect 112622 467004 112628 467016
rect 112487 466976 112628 467004
rect 112487 466973 112499 466976
rect 112441 466967 112499 466973
rect 112180 466936 112208 466967
rect 112622 466964 112628 466976
rect 112680 466964 112686 467016
rect 112806 466936 112812 466948
rect 112180 466908 112812 466936
rect 112806 466896 112812 466908
rect 112864 466896 112870 466948
rect 195054 466945 195060 466948
rect 195048 466899 195060 466945
rect 195112 466936 195118 466948
rect 195112 466908 195148 466936
rect 195054 466896 195060 466899
rect 195112 466896 195118 466908
rect 196161 466871 196219 466877
rect 196161 466837 196173 466871
rect 196207 466868 196219 466871
rect 340874 466868 340880 466880
rect 196207 466840 340880 466868
rect 196207 466837 196219 466840
rect 196161 466831 196219 466837
rect 340874 466828 340880 466840
rect 340932 466828 340938 466880
rect 207198 465400 207204 465452
rect 207256 465440 207262 465452
rect 223025 465443 223083 465449
rect 223025 465440 223037 465443
rect 207256 465412 223037 465440
rect 207256 465400 207262 465412
rect 223025 465409 223037 465412
rect 223071 465409 223083 465443
rect 223025 465403 223083 465409
rect 223117 465375 223175 465381
rect 223117 465341 223129 465375
rect 223163 465341 223175 465375
rect 223117 465335 223175 465341
rect 223301 465375 223359 465381
rect 223301 465341 223313 465375
rect 223347 465372 223359 465375
rect 223853 465375 223911 465381
rect 223853 465372 223865 465375
rect 223347 465344 223865 465372
rect 223347 465341 223359 465344
rect 223301 465335 223359 465341
rect 223853 465341 223865 465344
rect 223899 465341 223911 465375
rect 224402 465372 224408 465384
rect 224363 465344 224408 465372
rect 223853 465335 223911 465341
rect 120074 465196 120080 465248
rect 120132 465236 120138 465248
rect 222657 465239 222715 465245
rect 222657 465236 222669 465239
rect 120132 465208 222669 465236
rect 120132 465196 120138 465208
rect 222657 465205 222669 465208
rect 222703 465205 222715 465239
rect 223132 465236 223160 465335
rect 224402 465332 224408 465344
rect 224460 465372 224466 465384
rect 224460 465344 229094 465372
rect 224460 465332 224466 465344
rect 229066 465304 229094 465344
rect 255590 465304 255596 465316
rect 229066 465276 255596 465304
rect 255590 465264 255596 465276
rect 255648 465264 255654 465316
rect 311894 465236 311900 465248
rect 223132 465208 311900 465236
rect 222657 465199 222715 465205
rect 311894 465196 311900 465208
rect 311952 465196 311958 465248
rect 338022 463700 338028 463752
rect 338080 463740 338086 463752
rect 362773 463743 362831 463749
rect 362773 463740 362785 463743
rect 338080 463712 362785 463740
rect 338080 463700 338086 463712
rect 362773 463709 362785 463712
rect 362819 463709 362831 463743
rect 362773 463703 362831 463709
rect 6546 463020 6552 463072
rect 6604 463060 6610 463072
rect 109773 463063 109831 463069
rect 109773 463060 109785 463063
rect 6604 463032 109785 463060
rect 6604 463020 6610 463032
rect 109773 463029 109785 463032
rect 109819 463029 109831 463063
rect 109773 463023 109831 463029
rect 161446 460992 171134 461020
rect 3326 460912 3332 460964
rect 3384 460952 3390 460964
rect 161446 460952 161474 460992
rect 170398 460952 170404 460964
rect 3384 460924 161474 460952
rect 170359 460924 170404 460952
rect 3384 460912 3390 460924
rect 170398 460912 170404 460924
rect 170456 460912 170462 460964
rect 171106 460952 171134 460992
rect 358078 460952 358084 460964
rect 171106 460924 358084 460952
rect 358078 460912 358084 460924
rect 358136 460912 358142 460964
rect 185581 457623 185639 457629
rect 185581 457589 185593 457623
rect 185627 457620 185639 457623
rect 356698 457620 356704 457632
rect 185627 457592 356704 457620
rect 185627 457589 185639 457592
rect 185581 457583 185639 457589
rect 356698 457580 356704 457592
rect 356756 457580 356762 457632
rect 254210 457212 254216 457224
rect 254171 457184 254216 457212
rect 254210 457172 254216 457184
rect 254268 457172 254274 457224
rect 254118 457076 254124 457088
rect 254079 457048 254124 457076
rect 254118 457036 254124 457048
rect 254176 457036 254182 457088
rect 484210 455404 484216 455456
rect 484268 455444 484274 455456
rect 495434 455444 495440 455456
rect 484268 455416 495440 455444
rect 484268 455404 484274 455416
rect 495434 455404 495440 455416
rect 495492 455404 495498 455456
rect 133785 454359 133843 454365
rect 133785 454325 133797 454359
rect 133831 454356 133843 454359
rect 314286 454356 314292 454368
rect 133831 454328 314292 454356
rect 133831 454325 133843 454328
rect 133785 454319 133843 454325
rect 314286 454316 314292 454328
rect 314344 454316 314350 454368
rect 315298 453268 315304 453280
rect 315259 453240 315304 453268
rect 315298 453228 315304 453240
rect 315356 453228 315362 453280
rect 333514 451364 333520 451376
rect 45526 451336 53788 451364
rect 43162 451256 43168 451308
rect 43220 451296 43226 451308
rect 45526 451296 45554 451336
rect 53760 451305 53788 451336
rect 53852 451336 333520 451364
rect 43220 451268 45554 451296
rect 53635 451299 53693 451305
rect 43220 451256 43226 451268
rect 53635 451265 53647 451299
rect 53681 451296 53693 451299
rect 53745 451299 53803 451305
rect 53681 451265 53696 451296
rect 53635 451259 53696 451265
rect 53745 451265 53757 451299
rect 53791 451265 53803 451299
rect 53745 451259 53803 451265
rect 53668 451228 53696 451259
rect 53852 451228 53880 451336
rect 333514 451324 333520 451336
rect 333572 451324 333578 451376
rect 54018 451296 54024 451308
rect 53979 451268 54024 451296
rect 54018 451256 54024 451268
rect 54076 451256 54082 451308
rect 53668 451200 53880 451228
rect 53466 451092 53472 451104
rect 53427 451064 53472 451092
rect 53466 451052 53472 451064
rect 53524 451052 53530 451104
rect 53926 451092 53932 451104
rect 53887 451064 53932 451092
rect 53926 451052 53932 451064
rect 53984 451052 53990 451104
rect 142338 448536 142344 448588
rect 142396 448576 142402 448588
rect 175921 448579 175979 448585
rect 175921 448576 175933 448579
rect 142396 448548 175933 448576
rect 142396 448536 142402 448548
rect 175921 448545 175933 448548
rect 175967 448545 175979 448579
rect 175921 448539 175979 448545
rect 175734 448468 175740 448520
rect 175792 448517 175798 448520
rect 175792 448511 175841 448517
rect 175792 448477 175795 448511
rect 175829 448477 175841 448511
rect 176010 448508 176016 448520
rect 175971 448480 176016 448508
rect 175792 448471 175841 448477
rect 175792 448468 175798 448471
rect 176010 448468 176016 448480
rect 176068 448508 176074 448520
rect 419350 448508 419356 448520
rect 176068 448480 419356 448508
rect 176068 448468 176074 448480
rect 419350 448468 419356 448480
rect 419408 448468 419414 448520
rect 175550 448440 175556 448452
rect 175511 448412 175556 448440
rect 175550 448400 175556 448412
rect 175608 448400 175614 448452
rect 175642 448400 175648 448452
rect 175700 448440 175706 448452
rect 176197 448443 176255 448449
rect 175700 448412 175745 448440
rect 175700 448400 175706 448412
rect 176197 448409 176209 448443
rect 176243 448440 176255 448443
rect 178310 448440 178316 448452
rect 176243 448412 178316 448440
rect 176243 448409 176255 448412
rect 176197 448403 176255 448409
rect 178310 448400 178316 448412
rect 178368 448400 178374 448452
rect 175568 448372 175596 448400
rect 383838 448372 383844 448384
rect 175568 448344 383844 448372
rect 383838 448332 383844 448344
rect 383896 448332 383902 448384
rect 64782 447828 64788 447840
rect 64743 447800 64788 447828
rect 64782 447788 64788 447800
rect 64840 447788 64846 447840
rect 103486 446984 113174 447012
rect 53466 446904 53472 446956
rect 53524 446944 53530 446956
rect 103486 446944 103514 446984
rect 112254 446944 112260 446956
rect 53524 446916 103514 446944
rect 112215 446916 112260 446944
rect 53524 446904 53530 446916
rect 112254 446904 112260 446916
rect 112312 446904 112318 446956
rect 112346 446904 112352 446956
rect 112404 446944 112410 446956
rect 113146 446944 113174 446984
rect 334630 446947 334688 446953
rect 334630 446944 334642 446947
rect 112404 446916 112449 446944
rect 113146 446916 334642 446944
rect 112404 446904 112410 446916
rect 334630 446913 334642 446916
rect 334676 446913 334688 446947
rect 334630 446907 334688 446913
rect 112438 446876 112444 446888
rect 112399 446848 112444 446876
rect 112438 446836 112444 446848
rect 112496 446876 112502 446888
rect 140774 446876 140780 446888
rect 112496 446848 140780 446876
rect 112496 446836 112502 446848
rect 140774 446836 140780 446848
rect 140832 446836 140838 446888
rect 334897 446879 334955 446885
rect 334897 446845 334909 446879
rect 334943 446876 334955 446879
rect 383930 446876 383936 446888
rect 334943 446848 383936 446876
rect 334943 446845 334955 446848
rect 334897 446839 334955 446845
rect 383930 446836 383936 446848
rect 383988 446836 383994 446888
rect 88334 446700 88340 446752
rect 88392 446740 88398 446752
rect 111889 446743 111947 446749
rect 111889 446740 111901 446743
rect 88392 446712 111901 446740
rect 88392 446700 88398 446712
rect 111889 446709 111901 446712
rect 111935 446709 111947 446743
rect 333514 446740 333520 446752
rect 333475 446712 333520 446740
rect 111889 446703 111947 446709
rect 333514 446700 333520 446712
rect 333572 446700 333578 446752
rect 152366 443680 152372 443692
rect 152327 443652 152372 443680
rect 152366 443640 152372 443652
rect 152424 443640 152430 443692
rect 423858 443640 423864 443692
rect 423916 443680 423922 443692
rect 423953 443683 424011 443689
rect 423953 443680 423965 443683
rect 423916 443652 423965 443680
rect 423916 443640 423922 443652
rect 423953 443649 423965 443652
rect 423999 443649 424011 443683
rect 423953 443643 424011 443649
rect 152458 443612 152464 443624
rect 152419 443584 152464 443612
rect 152458 443572 152464 443584
rect 152516 443572 152522 443624
rect 152645 443615 152703 443621
rect 152645 443581 152657 443615
rect 152691 443612 152703 443615
rect 153197 443615 153255 443621
rect 153197 443612 153209 443615
rect 152691 443584 153209 443612
rect 152691 443581 152703 443584
rect 152645 443575 152703 443581
rect 153197 443581 153209 443584
rect 153243 443581 153255 443615
rect 153197 443575 153255 443581
rect 153841 443615 153899 443621
rect 153841 443581 153853 443615
rect 153887 443612 153899 443615
rect 154025 443615 154083 443621
rect 154025 443612 154037 443615
rect 153887 443584 154037 443612
rect 153887 443581 153899 443584
rect 153841 443575 153899 443581
rect 154025 443581 154037 443584
rect 154071 443612 154083 443615
rect 224402 443612 224408 443624
rect 154071 443584 224408 443612
rect 154071 443581 154083 443584
rect 154025 443575 154083 443581
rect 224402 443572 224408 443584
rect 224460 443572 224466 443624
rect 112622 443436 112628 443488
rect 112680 443476 112686 443488
rect 152001 443479 152059 443485
rect 152001 443476 152013 443479
rect 112680 443448 152013 443476
rect 112680 443436 112686 443448
rect 152001 443445 152013 443448
rect 152047 443445 152059 443479
rect 424042 443476 424048 443488
rect 424003 443448 424048 443476
rect 152001 443439 152059 443445
rect 424042 443436 424048 443448
rect 424100 443436 424106 443488
rect 152274 443096 152280 443148
rect 152332 443136 152338 443148
rect 152461 443139 152519 443145
rect 152461 443136 152473 443139
rect 152332 443108 152473 443136
rect 152332 443096 152338 443108
rect 152461 443105 152473 443108
rect 152507 443136 152519 443139
rect 154025 443139 154083 443145
rect 154025 443136 154037 443139
rect 152507 443108 154037 443136
rect 152507 443105 152519 443108
rect 152461 443099 152519 443105
rect 154025 443105 154037 443108
rect 154071 443105 154083 443139
rect 154025 443099 154083 443105
rect 153010 443000 153016 443012
rect 152971 442972 153016 443000
rect 153010 442960 153016 442972
rect 153068 442960 153074 443012
rect 281350 442592 281356 442604
rect 281311 442564 281356 442592
rect 281350 442552 281356 442564
rect 281408 442552 281414 442604
rect 376202 441980 376208 441992
rect 376163 441952 376208 441980
rect 376202 441940 376208 441952
rect 376260 441940 376266 441992
rect 376110 441844 376116 441856
rect 376071 441816 376116 441844
rect 376110 441804 376116 441816
rect 376168 441804 376174 441856
rect 311342 441600 311348 441652
rect 311400 441640 311406 441652
rect 495434 441640 495440 441652
rect 311400 441612 495440 441640
rect 311400 441600 311406 441612
rect 495434 441600 495440 441612
rect 495492 441600 495498 441652
rect 412082 439832 412088 439884
rect 412140 439872 412146 439884
rect 418525 439875 418583 439881
rect 418525 439872 418537 439875
rect 412140 439844 418537 439872
rect 412140 439832 412146 439844
rect 418525 439841 418537 439844
rect 418571 439841 418583 439875
rect 418525 439835 418583 439841
rect 42153 439807 42211 439813
rect 42153 439773 42165 439807
rect 42199 439804 42211 439807
rect 42429 439807 42487 439813
rect 42429 439804 42441 439807
rect 42199 439776 42441 439804
rect 42199 439773 42211 439776
rect 42153 439767 42211 439773
rect 42429 439773 42441 439776
rect 42475 439773 42487 439807
rect 42429 439767 42487 439773
rect 336550 439764 336556 439816
rect 336608 439804 336614 439816
rect 418433 439807 418491 439813
rect 418433 439804 418445 439807
rect 336608 439776 418445 439804
rect 336608 439764 336614 439776
rect 418433 439773 418445 439776
rect 418479 439773 418491 439807
rect 418433 439767 418491 439773
rect 418709 439807 418767 439813
rect 418709 439773 418721 439807
rect 418755 439773 418767 439807
rect 418709 439767 418767 439773
rect 43625 439739 43683 439745
rect 43625 439705 43637 439739
rect 43671 439736 43683 439739
rect 43993 439739 44051 439745
rect 43993 439736 44005 439739
rect 43671 439708 44005 439736
rect 43671 439705 43683 439708
rect 43625 439699 43683 439705
rect 43993 439705 44005 439708
rect 44039 439736 44051 439739
rect 195238 439736 195244 439748
rect 44039 439708 195244 439736
rect 44039 439705 44051 439708
rect 43993 439699 44051 439705
rect 195238 439696 195244 439708
rect 195296 439696 195302 439748
rect 412266 439696 412272 439748
rect 412324 439736 412330 439748
rect 418724 439736 418752 439767
rect 418798 439764 418804 439816
rect 418856 439804 418862 439816
rect 418856 439776 418901 439804
rect 418856 439764 418862 439776
rect 412324 439708 418752 439736
rect 412324 439696 412330 439708
rect 418982 439668 418988 439680
rect 418943 439640 418988 439668
rect 418982 439628 418988 439640
rect 419040 439628 419046 439680
rect 41969 439467 42027 439473
rect 41969 439433 41981 439467
rect 42015 439464 42027 439467
rect 42153 439467 42211 439473
rect 42153 439464 42165 439467
rect 42015 439436 42165 439464
rect 42015 439433 42027 439436
rect 41969 439427 42027 439433
rect 42153 439433 42165 439436
rect 42199 439433 42211 439467
rect 42153 439427 42211 439433
rect 43073 439467 43131 439473
rect 43073 439433 43085 439467
rect 43119 439464 43131 439467
rect 43162 439464 43168 439476
rect 43119 439436 43168 439464
rect 43119 439433 43131 439436
rect 43073 439427 43131 439433
rect 43162 439424 43168 439436
rect 43220 439424 43226 439476
rect 41782 439328 41788 439340
rect 41743 439300 41788 439328
rect 41782 439288 41788 439300
rect 41840 439288 41846 439340
rect 42521 439331 42579 439337
rect 42521 439297 42533 439331
rect 42567 439328 42579 439331
rect 43993 439331 44051 439337
rect 43993 439328 44005 439331
rect 42567 439300 44005 439328
rect 42567 439297 42579 439300
rect 42521 439291 42579 439297
rect 43993 439297 44005 439300
rect 44039 439297 44051 439331
rect 43993 439291 44051 439297
rect 281442 436908 281448 436960
rect 281500 436948 281506 436960
rect 397089 436951 397147 436957
rect 397089 436948 397101 436951
rect 281500 436920 397101 436948
rect 281500 436908 281506 436920
rect 397089 436917 397101 436920
rect 397135 436917 397147 436951
rect 397089 436911 397147 436917
rect 420638 435112 420644 435124
rect 47688 435084 420644 435112
rect 47688 435056 47716 435084
rect 420638 435072 420644 435084
rect 420696 435072 420702 435124
rect 47670 435044 47676 435056
rect 47583 435016 47676 435044
rect 47670 435004 47676 435016
rect 47728 435004 47734 435056
rect 47872 435016 56824 435044
rect 47688 434976 47716 435004
rect 47759 434979 47817 434985
rect 47759 434976 47771 434979
rect 47688 434948 47771 434976
rect 47759 434945 47771 434948
rect 47805 434945 47817 434979
rect 47759 434939 47817 434945
rect 44082 434868 44088 434920
rect 44140 434908 44146 434920
rect 47872 434908 47900 435016
rect 48038 434976 48044 434988
rect 47999 434948 48044 434976
rect 48038 434936 48044 434948
rect 48096 434936 48102 434988
rect 48222 434976 48228 434988
rect 48183 434948 48228 434976
rect 48222 434936 48228 434948
rect 48280 434936 48286 434988
rect 56796 434985 56824 435016
rect 56781 434979 56839 434985
rect 56781 434945 56793 434979
rect 56827 434945 56839 434979
rect 56781 434939 56839 434945
rect 44140 434880 47900 434908
rect 44140 434868 44146 434880
rect 48130 434868 48136 434920
rect 48188 434908 48194 434920
rect 143074 434908 143080 434920
rect 48188 434880 143080 434908
rect 48188 434868 48194 434880
rect 143074 434868 143080 434880
rect 143132 434868 143138 434920
rect 47854 434840 47860 434852
rect 47815 434812 47860 434840
rect 47854 434800 47860 434812
rect 47912 434800 47918 434852
rect 47949 434843 48007 434849
rect 47949 434809 47961 434843
rect 47995 434840 48007 434843
rect 263686 434840 263692 434852
rect 47995 434812 263692 434840
rect 47995 434809 48007 434812
rect 47949 434803 48007 434809
rect 263686 434800 263692 434812
rect 263744 434800 263750 434852
rect 47581 434775 47639 434781
rect 47581 434741 47593 434775
rect 47627 434772 47639 434775
rect 436738 434772 436744 434784
rect 47627 434744 436744 434772
rect 47627 434741 47639 434744
rect 47581 434735 47639 434741
rect 436738 434732 436744 434744
rect 436796 434732 436802 434784
rect 91462 434296 91468 434308
rect 91423 434268 91468 434296
rect 91462 434256 91468 434268
rect 91520 434256 91526 434308
rect 91649 434299 91707 434305
rect 91649 434265 91661 434299
rect 91695 434265 91707 434299
rect 91649 434259 91707 434265
rect 91833 434299 91891 434305
rect 91833 434265 91845 434299
rect 91879 434296 91891 434299
rect 293678 434296 293684 434308
rect 91879 434268 293684 434296
rect 91879 434265 91891 434268
rect 91833 434259 91891 434265
rect 91664 434228 91692 434259
rect 293678 434256 293684 434268
rect 293736 434256 293742 434308
rect 159082 434228 159088 434240
rect 91664 434200 159088 434228
rect 159082 434188 159088 434200
rect 159140 434188 159146 434240
rect 64049 433415 64107 433421
rect 64049 433381 64061 433415
rect 64095 433412 64107 433415
rect 267734 433412 267740 433424
rect 64095 433384 267740 433412
rect 64095 433381 64107 433384
rect 64049 433375 64107 433381
rect 267734 433372 267740 433384
rect 267792 433372 267798 433424
rect 3326 433304 3332 433356
rect 3384 433344 3390 433356
rect 338758 433344 338764 433356
rect 3384 433316 338764 433344
rect 3384 433304 3390 433316
rect 338758 433304 338764 433316
rect 338816 433304 338822 433356
rect 281350 432188 281356 432200
rect 281263 432160 281356 432188
rect 281350 432148 281356 432160
rect 281408 432188 281414 432200
rect 308306 432188 308312 432200
rect 281408 432160 308312 432188
rect 281408 432148 281414 432160
rect 308306 432148 308312 432160
rect 308364 432148 308370 432200
rect 281626 432129 281632 432132
rect 281620 432083 281632 432129
rect 281684 432120 281690 432132
rect 281684 432092 281720 432120
rect 281626 432080 281632 432083
rect 281684 432080 281690 432092
rect 282730 432052 282736 432064
rect 282643 432024 282736 432052
rect 282730 432012 282736 432024
rect 282788 432052 282794 432064
rect 496538 432052 496544 432064
rect 282788 432024 496544 432052
rect 282788 432012 282794 432024
rect 496538 432012 496544 432024
rect 496596 432012 496602 432064
rect 133690 429496 133696 429548
rect 133748 429536 133754 429548
rect 142249 429539 142307 429545
rect 142249 429536 142261 429539
rect 133748 429508 142261 429536
rect 133748 429496 133754 429508
rect 142249 429505 142261 429508
rect 142295 429505 142307 429539
rect 142430 429536 142436 429548
rect 142391 429508 142436 429536
rect 142249 429499 142307 429505
rect 142430 429496 142436 429508
rect 142488 429496 142494 429548
rect 142338 429400 142344 429412
rect 142299 429372 142344 429400
rect 142338 429360 142344 429372
rect 142396 429360 142402 429412
rect 412266 428448 412272 428460
rect 412227 428420 412272 428448
rect 412266 428408 412272 428420
rect 412324 428408 412330 428460
rect 412358 428408 412364 428460
rect 412416 428448 412422 428460
rect 412416 428420 412461 428448
rect 412416 428408 412422 428420
rect 289998 428340 290004 428392
rect 290056 428380 290062 428392
rect 411993 428383 412051 428389
rect 411993 428380 412005 428383
rect 290056 428352 412005 428380
rect 290056 428340 290062 428352
rect 411993 428349 412005 428352
rect 412039 428349 412051 428383
rect 411993 428343 412051 428349
rect 412545 428315 412603 428321
rect 412545 428312 412557 428315
rect 393286 428284 412557 428312
rect 184566 428204 184572 428256
rect 184624 428244 184630 428256
rect 393286 428244 393314 428284
rect 412545 428281 412557 428284
rect 412591 428281 412603 428315
rect 412545 428275 412603 428281
rect 412082 428244 412088 428256
rect 184624 428216 393314 428244
rect 412043 428216 412088 428244
rect 184624 428204 184630 428216
rect 412082 428204 412088 428216
rect 412140 428204 412146 428256
rect 311802 426708 311808 426760
rect 311860 426748 311866 426760
rect 450541 426751 450599 426757
rect 450541 426748 450553 426751
rect 311860 426720 450553 426748
rect 311860 426708 311866 426720
rect 450541 426717 450553 426720
rect 450587 426717 450599 426751
rect 450541 426711 450599 426717
rect 3326 425144 3332 425196
rect 3384 425184 3390 425196
rect 6638 425184 6644 425196
rect 3384 425156 6644 425184
rect 3384 425144 3390 425156
rect 6638 425144 6644 425156
rect 6696 425144 6702 425196
rect 91462 425076 91468 425128
rect 91520 425116 91526 425128
rect 92382 425116 92388 425128
rect 91520 425088 92388 425116
rect 91520 425076 91526 425088
rect 92382 425076 92388 425088
rect 92440 425116 92446 425128
rect 95878 425116 95884 425128
rect 92440 425088 95884 425116
rect 92440 425076 92446 425088
rect 95878 425076 95884 425088
rect 95936 425076 95942 425128
rect 239140 424612 248414 424640
rect 239030 424532 239036 424584
rect 239088 424572 239094 424584
rect 239140 424581 239168 424612
rect 239125 424575 239183 424581
rect 239125 424572 239137 424575
rect 239088 424544 239137 424572
rect 239088 424532 239094 424544
rect 239125 424541 239137 424544
rect 239171 424541 239183 424575
rect 239125 424535 239183 424541
rect 239309 424575 239367 424581
rect 239309 424541 239321 424575
rect 239355 424541 239367 424575
rect 248386 424572 248414 424612
rect 449894 424572 449900 424584
rect 248386 424544 449900 424572
rect 239309 424535 239367 424541
rect 46014 424464 46020 424516
rect 46072 424504 46078 424516
rect 238941 424507 238999 424513
rect 238941 424504 238953 424507
rect 46072 424476 238953 424504
rect 46072 424464 46078 424476
rect 238941 424473 238953 424476
rect 238987 424473 238999 424507
rect 239324 424504 239352 424535
rect 449894 424532 449900 424544
rect 449952 424532 449958 424584
rect 312078 424504 312084 424516
rect 239324 424476 312084 424504
rect 238941 424467 238999 424473
rect 312078 424464 312084 424476
rect 312136 424464 312142 424516
rect 312078 423648 312084 423700
rect 312136 423688 312142 423700
rect 495986 423688 495992 423700
rect 312136 423660 495992 423688
rect 312136 423648 312142 423660
rect 495986 423648 495992 423660
rect 496044 423648 496050 423700
rect 15010 423512 15016 423564
rect 15068 423552 15074 423564
rect 331398 423552 331404 423564
rect 15068 423524 316034 423552
rect 331311 423524 331404 423552
rect 15068 423512 15074 423524
rect 132586 423444 132592 423496
rect 132644 423484 132650 423496
rect 133690 423484 133696 423496
rect 132644 423456 133696 423484
rect 132644 423444 132650 423456
rect 133690 423444 133696 423456
rect 133748 423444 133754 423496
rect 133874 423484 133880 423496
rect 133835 423456 133880 423484
rect 133874 423444 133880 423456
rect 133932 423444 133938 423496
rect 133966 423444 133972 423496
rect 134024 423484 134030 423496
rect 134150 423493 134156 423496
rect 134107 423487 134156 423493
rect 134024 423456 134069 423484
rect 134024 423444 134030 423456
rect 134107 423453 134119 423487
rect 134153 423453 134156 423487
rect 134107 423447 134156 423453
rect 134150 423444 134156 423447
rect 134208 423444 134214 423496
rect 134245 423487 134303 423493
rect 134245 423453 134257 423487
rect 134291 423484 134303 423487
rect 316006 423484 316034 423524
rect 331398 423512 331404 423524
rect 331456 423552 331462 423564
rect 332045 423555 332103 423561
rect 332045 423552 332057 423555
rect 331456 423524 332057 423552
rect 331456 423512 331462 423524
rect 332045 423521 332057 423524
rect 332091 423521 332103 423555
rect 332045 423515 332103 423521
rect 331125 423487 331183 423493
rect 331125 423484 331137 423487
rect 134291 423456 142154 423484
rect 316006 423456 331137 423484
rect 134291 423453 134303 423456
rect 134245 423447 134303 423453
rect 142126 423416 142154 423456
rect 331125 423453 331137 423456
rect 331171 423453 331183 423487
rect 331125 423447 331183 423453
rect 331214 423444 331220 423496
rect 331272 423484 331278 423496
rect 331308 423487 331366 423493
rect 331308 423484 331320 423487
rect 331272 423456 331320 423484
rect 331272 423444 331278 423456
rect 331308 423453 331320 423456
rect 331354 423453 331366 423487
rect 331308 423447 331366 423453
rect 331490 423444 331496 423496
rect 331548 423484 331554 423496
rect 331548 423456 331593 423484
rect 331548 423444 331554 423456
rect 331674 423444 331680 423496
rect 331732 423484 331738 423496
rect 331732 423456 335354 423484
rect 331732 423444 331738 423456
rect 244458 423416 244464 423428
rect 122806 423388 137324 423416
rect 142126 423388 244464 423416
rect 89254 423308 89260 423360
rect 89312 423348 89318 423360
rect 122806 423348 122834 423388
rect 134334 423348 134340 423360
rect 89312 423320 122834 423348
rect 134295 423320 134340 423348
rect 89312 423308 89318 423320
rect 134334 423308 134340 423320
rect 134392 423308 134398 423360
rect 137296 423348 137324 423388
rect 244458 423376 244464 423388
rect 244516 423376 244522 423428
rect 335326 423416 335354 423456
rect 385126 423416 385132 423428
rect 335326 423388 385132 423416
rect 385126 423376 385132 423388
rect 385184 423376 385190 423428
rect 331769 423351 331827 423357
rect 331769 423348 331781 423351
rect 137296 423320 331781 423348
rect 331769 423317 331781 423320
rect 331815 423317 331827 423351
rect 331769 423311 331827 423317
rect 27522 423144 27528 423156
rect 27483 423116 27528 423144
rect 27522 423104 27528 423116
rect 27580 423104 27586 423156
rect 133966 423104 133972 423156
rect 134024 423144 134030 423156
rect 205266 423144 205272 423156
rect 134024 423116 205272 423144
rect 134024 423104 134030 423116
rect 205266 423104 205272 423116
rect 205324 423104 205330 423156
rect 332045 423147 332103 423153
rect 332045 423113 332057 423147
rect 332091 423144 332103 423147
rect 451458 423144 451464 423156
rect 332091 423116 451464 423144
rect 332091 423113 332103 423116
rect 332045 423107 332103 423113
rect 451458 423104 451464 423116
rect 451516 423104 451522 423156
rect 32033 423079 32091 423085
rect 32033 423076 32045 423079
rect 27448 423048 32045 423076
rect 27448 423020 27476 423048
rect 32033 423045 32045 423048
rect 32079 423045 32091 423079
rect 32033 423039 32091 423045
rect 134150 423036 134156 423088
rect 134208 423076 134214 423088
rect 205358 423076 205364 423088
rect 134208 423048 205364 423076
rect 134208 423036 134214 423048
rect 205358 423036 205364 423048
rect 205416 423036 205422 423088
rect 27430 423008 27436 423020
rect 27391 422980 27436 423008
rect 27430 422968 27436 422980
rect 27488 422968 27494 423020
rect 27985 423011 28043 423017
rect 27985 422977 27997 423011
rect 28031 422977 28043 423011
rect 27985 422971 28043 422977
rect 28261 423011 28319 423017
rect 28261 422977 28273 423011
rect 28307 423008 28319 423011
rect 92382 423008 92388 423020
rect 28307 422980 92388 423008
rect 28307 422977 28319 422980
rect 28261 422971 28319 422977
rect 27617 422943 27675 422949
rect 27617 422909 27629 422943
rect 27663 422909 27675 422943
rect 28000 422940 28028 422971
rect 92382 422968 92388 422980
rect 92440 422968 92446 423020
rect 28353 422943 28411 422949
rect 28353 422940 28365 422943
rect 28000 422912 28365 422940
rect 27617 422903 27675 422909
rect 28353 422909 28365 422912
rect 28399 422909 28411 422943
rect 120994 422940 121000 422952
rect 28353 422903 28411 422909
rect 31772 422912 121000 422940
rect 27632 422872 27660 422903
rect 31772 422872 31800 422912
rect 120994 422900 121000 422912
rect 121052 422900 121058 422952
rect 67358 422872 67364 422884
rect 27632 422844 31800 422872
rect 31956 422844 67364 422872
rect 28353 422807 28411 422813
rect 28353 422773 28365 422807
rect 28399 422804 28411 422807
rect 31956 422804 31984 422844
rect 67358 422832 67364 422844
rect 67416 422832 67422 422884
rect 28399 422776 31984 422804
rect 32033 422807 32091 422813
rect 28399 422773 28411 422776
rect 28353 422767 28411 422773
rect 32033 422773 32045 422807
rect 32079 422804 32091 422807
rect 55398 422804 55404 422816
rect 32079 422776 55404 422804
rect 32079 422773 32091 422776
rect 32033 422767 32091 422773
rect 55398 422764 55404 422776
rect 55456 422764 55462 422816
rect 9674 422560 9680 422612
rect 9732 422600 9738 422612
rect 133874 422600 133880 422612
rect 9732 422572 133880 422600
rect 9732 422560 9738 422572
rect 133874 422560 133880 422572
rect 133932 422560 133938 422612
rect 443914 421308 443920 421320
rect 443827 421280 443920 421308
rect 443914 421268 443920 421280
rect 443972 421308 443978 421320
rect 470410 421308 470416 421320
rect 443972 421280 470416 421308
rect 443972 421268 443978 421280
rect 470410 421268 470416 421280
rect 470468 421268 470474 421320
rect 338206 421200 338212 421252
rect 338264 421240 338270 421252
rect 443650 421243 443708 421249
rect 443650 421240 443662 421243
rect 338264 421212 443662 421240
rect 338264 421200 338270 421212
rect 443650 421209 443662 421212
rect 443696 421209 443708 421243
rect 443650 421203 443708 421209
rect 442534 421172 442540 421184
rect 442495 421144 442540 421172
rect 442534 421132 442540 421144
rect 442592 421132 442598 421184
rect 3970 417528 3976 417580
rect 4028 417568 4034 417580
rect 333977 417571 334035 417577
rect 333977 417568 333989 417571
rect 4028 417540 333989 417568
rect 4028 417528 4034 417540
rect 333977 417537 333989 417540
rect 334023 417537 334035 417571
rect 333977 417531 334035 417537
rect 334066 417528 334072 417580
rect 334124 417568 334130 417580
rect 334124 417540 334169 417568
rect 334124 417528 334130 417540
rect 334342 417500 334348 417512
rect 334303 417472 334348 417500
rect 334342 417460 334348 417472
rect 334400 417460 334406 417512
rect 203058 417392 203064 417444
rect 203116 417432 203122 417444
rect 334253 417435 334311 417441
rect 334253 417432 334265 417435
rect 203116 417404 334265 417432
rect 203116 417392 203122 417404
rect 334253 417401 334265 417404
rect 334299 417401 334311 417435
rect 334253 417395 334311 417401
rect 5074 417324 5080 417376
rect 5132 417364 5138 417376
rect 333793 417367 333851 417373
rect 333793 417364 333805 417367
rect 5132 417336 333805 417364
rect 5132 417324 5138 417336
rect 333793 417333 333805 417336
rect 333839 417333 333851 417367
rect 333793 417327 333851 417333
rect 136542 417160 136548 417172
rect 136503 417132 136548 417160
rect 136542 417120 136548 417132
rect 136600 417120 136606 417172
rect 152458 415488 152464 415540
rect 152516 415528 152522 415540
rect 256513 415531 256571 415537
rect 256513 415528 256525 415531
rect 152516 415500 256525 415528
rect 152516 415488 152522 415500
rect 256513 415497 256525 415500
rect 256559 415497 256571 415531
rect 256513 415491 256571 415497
rect 101490 415420 101496 415472
rect 101548 415460 101554 415472
rect 256881 415463 256939 415469
rect 256881 415460 256893 415463
rect 101548 415432 256893 415460
rect 101548 415420 101554 415432
rect 256881 415429 256893 415432
rect 256927 415429 256939 415463
rect 279697 415463 279755 415469
rect 279697 415460 279709 415463
rect 256881 415423 256939 415429
rect 279528 415432 279709 415460
rect 279234 415392 279240 415404
rect 279195 415364 279240 415392
rect 279234 415352 279240 415364
rect 279292 415352 279298 415404
rect 279329 415395 279387 415401
rect 279329 415361 279341 415395
rect 279375 415392 279387 415395
rect 279528 415392 279556 415432
rect 279697 415429 279709 415432
rect 279743 415429 279755 415463
rect 346854 415460 346860 415472
rect 279697 415423 279755 415429
rect 279804 415432 346860 415460
rect 279375 415364 279556 415392
rect 279375 415361 279387 415364
rect 279329 415355 279387 415361
rect 8110 415284 8116 415336
rect 8168 415324 8174 415336
rect 256973 415327 257031 415333
rect 256973 415324 256985 415327
rect 8168 415296 256985 415324
rect 8168 415284 8174 415296
rect 256973 415293 256985 415296
rect 257019 415293 257031 415327
rect 256973 415287 257031 415293
rect 257062 415284 257068 415336
rect 257120 415324 257126 415336
rect 262490 415324 262496 415336
rect 257120 415296 262496 415324
rect 257120 415284 257126 415296
rect 262490 415284 262496 415296
rect 262548 415284 262554 415336
rect 279053 415327 279111 415333
rect 279053 415324 279065 415327
rect 267706 415296 279065 415324
rect 232130 415216 232136 415268
rect 232188 415256 232194 415268
rect 267706 415256 267734 415296
rect 279053 415293 279065 415296
rect 279099 415293 279111 415327
rect 279602 415324 279608 415336
rect 279515 415296 279608 415324
rect 279053 415287 279111 415293
rect 279602 415284 279608 415296
rect 279660 415324 279666 415336
rect 279804 415324 279832 415432
rect 346854 415420 346860 415432
rect 346912 415420 346918 415472
rect 279881 415395 279939 415401
rect 279881 415361 279893 415395
rect 279927 415392 279939 415395
rect 346578 415392 346584 415404
rect 279927 415364 346584 415392
rect 279927 415361 279939 415364
rect 279881 415355 279939 415361
rect 346578 415352 346584 415364
rect 346636 415352 346642 415404
rect 279660 415296 279832 415324
rect 279660 415284 279666 415296
rect 279513 415259 279571 415265
rect 279513 415256 279525 415259
rect 232188 415228 267734 415256
rect 277366 415228 279525 415256
rect 232188 415216 232194 415228
rect 95602 415148 95608 415200
rect 95660 415188 95666 415200
rect 277366 415188 277394 415228
rect 279513 415225 279525 415228
rect 279559 415225 279571 415259
rect 279513 415219 279571 415225
rect 95660 415160 277394 415188
rect 95660 415148 95666 415160
rect 119614 414780 119620 414792
rect 119575 414752 119620 414780
rect 119614 414740 119620 414752
rect 119672 414740 119678 414792
rect 318058 414264 318064 414316
rect 318116 414304 318122 414316
rect 402681 414307 402739 414313
rect 402681 414304 402693 414307
rect 318116 414276 402693 414304
rect 318116 414264 318122 414276
rect 402681 414273 402693 414276
rect 402727 414273 402739 414307
rect 402681 414267 402739 414273
rect 402422 414236 402428 414248
rect 402383 414208 402428 414236
rect 402422 414196 402428 414208
rect 402480 414196 402486 414248
rect 403802 414100 403808 414112
rect 403715 414072 403808 414100
rect 403802 414060 403808 414072
rect 403860 414100 403866 414112
rect 485590 414100 485596 414112
rect 403860 414072 485596 414100
rect 403860 414060 403866 414072
rect 485590 414060 485596 414072
rect 485648 414060 485654 414112
rect 258902 413896 258908 413908
rect 258863 413868 258908 413896
rect 258902 413856 258908 413868
rect 258960 413856 258966 413908
rect 260285 413695 260343 413701
rect 260285 413661 260297 413695
rect 260331 413692 260343 413695
rect 281350 413692 281356 413704
rect 260331 413664 281356 413692
rect 260331 413661 260343 413664
rect 260285 413655 260343 413661
rect 281350 413652 281356 413664
rect 281408 413652 281414 413704
rect 205634 413584 205640 413636
rect 205692 413624 205698 413636
rect 260018 413627 260076 413633
rect 260018 413624 260030 413627
rect 205692 413596 260030 413624
rect 205692 413584 205698 413596
rect 260018 413593 260030 413596
rect 260064 413593 260076 413627
rect 260018 413587 260076 413593
rect 143810 412808 143816 412820
rect 143771 412780 143816 412808
rect 143810 412768 143816 412780
rect 143868 412768 143874 412820
rect 254118 412632 254124 412684
rect 254176 412672 254182 412684
rect 257430 412672 257436 412684
rect 254176 412644 257436 412672
rect 254176 412632 254182 412644
rect 257430 412632 257436 412644
rect 257488 412632 257494 412684
rect 151449 411927 151507 411933
rect 151449 411893 151461 411927
rect 151495 411924 151507 411927
rect 389174 411924 389180 411936
rect 151495 411896 389180 411924
rect 151495 411893 151507 411896
rect 151449 411887 151507 411893
rect 389174 411884 389180 411896
rect 389232 411884 389238 411936
rect 4062 411476 4068 411528
rect 4120 411516 4126 411528
rect 338393 411519 338451 411525
rect 338393 411516 338405 411519
rect 4120 411488 338405 411516
rect 4120 411476 4126 411488
rect 338393 411485 338405 411488
rect 338439 411485 338451 411519
rect 338393 411479 338451 411485
rect 99650 411040 99656 411052
rect 99611 411012 99656 411040
rect 99650 411000 99656 411012
rect 99708 411000 99714 411052
rect 99834 411040 99840 411052
rect 99795 411012 99840 411040
rect 99834 411000 99840 411012
rect 99892 411000 99898 411052
rect 99668 410972 99696 411000
rect 254118 410972 254124 410984
rect 99668 410944 254124 410972
rect 254118 410932 254124 410944
rect 254176 410932 254182 410984
rect 99929 410907 99987 410913
rect 99929 410873 99941 410907
rect 99975 410904 99987 410907
rect 325786 410904 325792 410916
rect 99975 410876 325792 410904
rect 99975 410873 99987 410876
rect 99929 410867 99987 410873
rect 112530 410632 112536 410644
rect 112491 410604 112536 410632
rect 112530 410592 112536 410604
rect 112588 410592 112594 410644
rect 112990 410632 112996 410644
rect 112951 410604 112996 410632
rect 112990 410592 112996 410604
rect 113048 410592 113054 410644
rect 325666 410632 325694 410876
rect 325786 410864 325792 410876
rect 325844 410864 325850 410916
rect 335538 410632 335544 410644
rect 325666 410604 335544 410632
rect 335538 410592 335544 410604
rect 335596 410592 335602 410644
rect 99834 410524 99840 410576
rect 99892 410564 99898 410576
rect 331490 410564 331496 410576
rect 99892 410536 331496 410564
rect 99892 410524 99898 410536
rect 331490 410524 331496 410536
rect 331548 410524 331554 410576
rect 113082 410496 113088 410508
rect 113043 410468 113088 410496
rect 113082 410456 113088 410468
rect 113140 410456 113146 410508
rect 112717 410431 112775 410437
rect 112717 410397 112729 410431
rect 112763 410397 112775 410431
rect 112717 410391 112775 410397
rect 112732 410360 112760 410391
rect 112806 410388 112812 410440
rect 112864 410428 112870 410440
rect 375374 410428 375380 410440
rect 112864 410400 112909 410428
rect 113146 410400 375380 410428
rect 112864 410388 112870 410400
rect 113146 410360 113174 410400
rect 375374 410388 375380 410400
rect 375432 410428 375438 410440
rect 375650 410428 375656 410440
rect 375432 410400 375656 410428
rect 375432 410388 375438 410400
rect 375650 410388 375656 410400
rect 375708 410388 375714 410440
rect 253106 410360 253112 410372
rect 112732 410332 113174 410360
rect 122806 410332 253112 410360
rect 112806 410252 112812 410304
rect 112864 410292 112870 410304
rect 122806 410292 122834 410332
rect 253106 410320 253112 410332
rect 253164 410320 253170 410372
rect 112864 410264 122834 410292
rect 112864 410252 112870 410264
rect 55508 409992 64874 410020
rect 55508 409964 55536 409992
rect 55306 409952 55312 409964
rect 55267 409924 55312 409952
rect 55306 409912 55312 409924
rect 55364 409912 55370 409964
rect 55490 409952 55496 409964
rect 55451 409924 55496 409952
rect 55490 409912 55496 409924
rect 55548 409912 55554 409964
rect 55677 409955 55735 409961
rect 55677 409921 55689 409955
rect 55723 409921 55735 409955
rect 64846 409952 64874 409992
rect 198458 409952 198464 409964
rect 64846 409924 198464 409952
rect 55677 409915 55735 409921
rect 55692 409884 55720 409915
rect 198458 409912 198464 409924
rect 198516 409912 198522 409964
rect 89438 409884 89444 409896
rect 55692 409856 89444 409884
rect 89438 409844 89444 409856
rect 89496 409844 89502 409896
rect 57793 409547 57851 409553
rect 57793 409544 57805 409547
rect 57256 409516 57805 409544
rect 57146 409408 57152 409420
rect 57107 409380 57152 409408
rect 57146 409368 57152 409380
rect 57204 409368 57210 409420
rect 57256 409417 57284 409516
rect 57793 409513 57805 409516
rect 57839 409513 57851 409547
rect 57793 409507 57851 409513
rect 57241 409411 57299 409417
rect 57241 409377 57253 409411
rect 57287 409377 57299 409411
rect 57241 409371 57299 409377
rect 57330 409368 57336 409420
rect 57388 409408 57394 409420
rect 342898 409408 342904 409420
rect 57388 409380 342904 409408
rect 57388 409368 57394 409380
rect 342898 409368 342904 409380
rect 342956 409368 342962 409420
rect 56870 409340 56876 409352
rect 56831 409312 56876 409340
rect 56870 409300 56876 409312
rect 56928 409300 56934 409352
rect 56965 409343 57023 409349
rect 56965 409309 56977 409343
rect 57011 409309 57023 409343
rect 177298 409340 177304 409352
rect 56965 409303 57023 409309
rect 57348 409312 177304 409340
rect 56686 409204 56692 409216
rect 56647 409176 56692 409204
rect 56686 409164 56692 409176
rect 56744 409164 56750 409216
rect 56980 409204 57008 409303
rect 57348 409204 57376 409312
rect 177298 409300 177304 409312
rect 177356 409300 177362 409352
rect 57793 409275 57851 409281
rect 57793 409241 57805 409275
rect 57839 409272 57851 409275
rect 92290 409272 92296 409284
rect 57839 409244 92296 409272
rect 57839 409241 57851 409244
rect 57793 409235 57851 409241
rect 92290 409232 92296 409244
rect 92348 409232 92354 409284
rect 90634 409204 90640 409216
rect 56980 409176 57376 409204
rect 64846 409176 90640 409204
rect 56870 408960 56876 409012
rect 56928 409000 56934 409012
rect 64846 409000 64874 409176
rect 90634 409164 90640 409176
rect 90692 409164 90698 409216
rect 56928 408972 64874 409000
rect 56928 408960 56934 408972
rect 3326 407124 3332 407176
rect 3384 407164 3390 407176
rect 11698 407164 11704 407176
rect 3384 407136 11704 407164
rect 3384 407124 3390 407136
rect 11698 407124 11704 407136
rect 11756 407124 11762 407176
rect 316862 407124 316868 407176
rect 316920 407164 316926 407176
rect 495434 407164 495440 407176
rect 316920 407136 495440 407164
rect 316920 407124 316926 407136
rect 495434 407124 495440 407136
rect 495492 407124 495498 407176
rect 3326 406988 3332 407040
rect 3384 407028 3390 407040
rect 4062 407028 4068 407040
rect 3384 407000 4068 407028
rect 3384 406988 3390 407000
rect 4062 406988 4068 407000
rect 4120 406988 4126 407040
rect 35802 406036 35808 406088
rect 35860 406076 35866 406088
rect 441801 406079 441859 406085
rect 441801 406076 441813 406079
rect 35860 406048 441813 406076
rect 35860 406036 35866 406048
rect 441801 406045 441813 406048
rect 441847 406045 441859 406079
rect 441801 406039 441859 406045
rect 114094 405600 114100 405612
rect 114055 405572 114100 405600
rect 114094 405560 114100 405572
rect 114152 405560 114158 405612
rect 3050 403180 3056 403232
rect 3108 403220 3114 403232
rect 56597 403223 56655 403229
rect 56597 403220 56609 403223
rect 3108 403192 56609 403220
rect 3108 403180 3114 403192
rect 56597 403189 56609 403192
rect 56643 403189 56655 403223
rect 56597 403183 56655 403189
rect 170398 402908 170404 402960
rect 170456 402948 170462 402960
rect 495434 402948 495440 402960
rect 170456 402920 495440 402948
rect 170456 402908 170462 402920
rect 495434 402908 495440 402920
rect 495492 402908 495498 402960
rect 119982 401684 119988 401736
rect 120040 401724 120046 401736
rect 169941 401727 169999 401733
rect 169941 401724 169953 401727
rect 120040 401696 169953 401724
rect 120040 401684 120046 401696
rect 169941 401693 169953 401696
rect 169987 401693 169999 401727
rect 169941 401687 169999 401693
rect 2958 401616 2964 401668
rect 3016 401656 3022 401668
rect 312170 401656 312176 401668
rect 3016 401628 312176 401656
rect 3016 401616 3022 401628
rect 312170 401616 312176 401628
rect 312228 401616 312234 401668
rect 67177 400707 67235 400713
rect 67177 400673 67189 400707
rect 67223 400704 67235 400707
rect 414290 400704 414296 400716
rect 67223 400676 414296 400704
rect 67223 400673 67235 400676
rect 67177 400667 67235 400673
rect 414290 400664 414296 400676
rect 414348 400664 414354 400716
rect 67082 400636 67088 400648
rect 67043 400608 67088 400636
rect 67082 400596 67088 400608
rect 67140 400596 67146 400648
rect 67358 400636 67364 400648
rect 67319 400608 67364 400636
rect 67358 400596 67364 400608
rect 67416 400596 67422 400648
rect 67450 400596 67456 400648
rect 67508 400636 67514 400648
rect 67508 400608 67553 400636
rect 67508 400596 67514 400608
rect 67634 400596 67640 400648
rect 67692 400636 67698 400648
rect 423766 400636 423772 400648
rect 67692 400608 423772 400636
rect 67692 400596 67698 400608
rect 423766 400596 423772 400608
rect 423824 400596 423830 400648
rect 67100 400568 67128 400596
rect 283282 400568 283288 400580
rect 67100 400540 283288 400568
rect 283282 400528 283288 400540
rect 283340 400528 283346 400580
rect 67634 400500 67640 400512
rect 67595 400472 67640 400500
rect 67634 400460 67640 400472
rect 67692 400460 67698 400512
rect 268933 399959 268991 399965
rect 268933 399925 268945 399959
rect 268979 399956 268991 399959
rect 314378 399956 314384 399968
rect 268979 399928 314384 399956
rect 268979 399925 268991 399928
rect 268933 399919 268991 399925
rect 314378 399916 314384 399928
rect 314436 399916 314442 399968
rect 252925 399551 252983 399557
rect 252925 399517 252937 399551
rect 252971 399548 252983 399551
rect 375466 399548 375472 399560
rect 252971 399520 375472 399548
rect 252971 399517 252983 399520
rect 252925 399511 252983 399517
rect 375466 399508 375472 399520
rect 375524 399548 375530 399560
rect 376110 399548 376116 399560
rect 375524 399520 376116 399548
rect 375524 399508 375530 399520
rect 376110 399508 376116 399520
rect 376168 399508 376174 399560
rect 253106 399412 253112 399424
rect 253019 399384 253112 399412
rect 253106 399372 253112 399384
rect 253164 399412 253170 399424
rect 426710 399412 426716 399424
rect 253164 399384 426716 399412
rect 253164 399372 253170 399384
rect 426710 399372 426716 399384
rect 426768 399372 426774 399424
rect 400030 398460 400036 398472
rect 399991 398432 400036 398460
rect 400030 398420 400036 398432
rect 400088 398420 400094 398472
rect 326522 397780 326528 397792
rect 326483 397752 326528 397780
rect 326522 397740 326528 397752
rect 326580 397740 326586 397792
rect 316954 397536 316960 397588
rect 317012 397576 317018 397588
rect 495434 397576 495440 397588
rect 317012 397548 495440 397576
rect 317012 397536 317018 397548
rect 495434 397536 495440 397548
rect 495492 397536 495498 397588
rect 211062 397468 211068 397520
rect 211120 397508 211126 397520
rect 340785 397511 340843 397517
rect 340785 397508 340797 397511
rect 211120 397480 340797 397508
rect 211120 397468 211126 397480
rect 340785 397477 340797 397480
rect 340831 397477 340843 397511
rect 340785 397471 340843 397477
rect 282641 396287 282699 396293
rect 282641 396253 282653 396287
rect 282687 396284 282699 396287
rect 398098 396284 398104 396296
rect 282687 396256 398104 396284
rect 282687 396253 282699 396256
rect 282641 396247 282699 396253
rect 398098 396244 398104 396256
rect 398156 396244 398162 396296
rect 43070 395808 43076 395820
rect 43031 395780 43076 395808
rect 43070 395768 43076 395780
rect 43128 395768 43134 395820
rect 3786 395564 3792 395616
rect 3844 395604 3850 395616
rect 313737 395607 313795 395613
rect 313737 395604 313749 395607
rect 3844 395576 313749 395604
rect 3844 395564 3850 395576
rect 313737 395573 313749 395576
rect 313783 395573 313795 395607
rect 313737 395567 313795 395573
rect 380529 395267 380587 395273
rect 380529 395233 380541 395267
rect 380575 395264 380587 395267
rect 380618 395264 380624 395276
rect 380575 395236 380624 395264
rect 380575 395233 380587 395236
rect 380529 395227 380587 395233
rect 380618 395224 380624 395236
rect 380676 395224 380682 395276
rect 11790 395196 11796 395208
rect 11751 395168 11796 395196
rect 11790 395156 11796 395168
rect 11848 395156 11854 395208
rect 380710 395196 380716 395208
rect 380671 395168 380716 395196
rect 380710 395156 380716 395168
rect 380768 395156 380774 395208
rect 373966 395100 383654 395128
rect 11977 395063 12035 395069
rect 11977 395029 11989 395063
rect 12023 395060 12035 395063
rect 373966 395060 373994 395100
rect 380894 395060 380900 395072
rect 12023 395032 373994 395060
rect 380855 395032 380900 395060
rect 12023 395029 12035 395032
rect 11977 395023 12035 395029
rect 380894 395020 380900 395032
rect 380952 395020 380958 395072
rect 383626 395060 383654 395100
rect 433978 395060 433984 395072
rect 383626 395032 433984 395060
rect 433978 395020 433984 395032
rect 434036 395020 434042 395072
rect 22830 394856 22836 394868
rect 22791 394828 22836 394856
rect 22830 394816 22836 394828
rect 22888 394856 22894 394868
rect 23385 394859 23443 394865
rect 23385 394856 23397 394859
rect 22888 394828 23397 394856
rect 22888 394816 22894 394828
rect 23385 394825 23397 394828
rect 23431 394825 23443 394859
rect 23385 394819 23443 394825
rect 45738 394788 45744 394800
rect 23032 394760 45744 394788
rect 22922 394680 22928 394732
rect 22980 394720 22986 394732
rect 23032 394729 23060 394760
rect 45738 394748 45744 394760
rect 45796 394748 45802 394800
rect 23017 394723 23075 394729
rect 23017 394720 23029 394723
rect 22980 394692 23029 394720
rect 22980 394680 22986 394692
rect 23017 394689 23029 394692
rect 23063 394689 23075 394723
rect 23017 394683 23075 394689
rect 23385 394723 23443 394729
rect 23385 394689 23397 394723
rect 23431 394720 23443 394723
rect 360378 394720 360384 394732
rect 23431 394692 360384 394720
rect 23431 394689 23443 394692
rect 23385 394683 23443 394689
rect 360378 394680 360384 394692
rect 360436 394680 360442 394732
rect 452102 394176 452108 394188
rect 452063 394148 452108 394176
rect 452102 394136 452108 394148
rect 452160 394136 452166 394188
rect 451918 394108 451924 394120
rect 451879 394080 451924 394108
rect 451918 394068 451924 394080
rect 451976 394068 451982 394120
rect 452013 394043 452071 394049
rect 452013 394040 452025 394043
rect 431926 394012 452025 394040
rect 167822 393728 167828 393780
rect 167880 393768 167886 393780
rect 431926 393768 431954 394012
rect 452013 394009 452025 394012
rect 452059 394009 452071 394043
rect 452013 394003 452071 394009
rect 451550 393972 451556 393984
rect 451511 393944 451556 393972
rect 451550 393932 451556 393944
rect 451608 393932 451614 393984
rect 167880 393740 431954 393768
rect 167880 393728 167886 393740
rect 6086 393388 6092 393440
rect 6144 393428 6150 393440
rect 20533 393431 20591 393437
rect 20533 393428 20545 393431
rect 6144 393400 20545 393428
rect 6144 393388 6150 393400
rect 20533 393397 20545 393400
rect 20579 393397 20591 393431
rect 20533 393391 20591 393397
rect 257065 392343 257123 392349
rect 257065 392309 257077 392343
rect 257111 392340 257123 392343
rect 330478 392340 330484 392352
rect 257111 392312 330484 392340
rect 257111 392309 257123 392312
rect 257065 392303 257123 392309
rect 330478 392300 330484 392312
rect 330536 392300 330542 392352
rect 3602 389648 3608 389700
rect 3660 389688 3666 389700
rect 3786 389688 3792 389700
rect 3660 389660 3792 389688
rect 3660 389648 3666 389660
rect 3786 389648 3792 389660
rect 3844 389648 3850 389700
rect 3602 389172 3608 389224
rect 3660 389212 3666 389224
rect 214558 389212 214564 389224
rect 3660 389184 214564 389212
rect 3660 389172 3666 389184
rect 214558 389172 214564 389184
rect 214616 389172 214622 389224
rect 346762 387648 346768 387660
rect 346723 387620 346768 387648
rect 346762 387608 346768 387620
rect 346820 387608 346826 387660
rect 346854 387608 346860 387660
rect 346912 387648 346918 387660
rect 346912 387620 354674 387648
rect 346912 387608 346918 387620
rect 346486 387580 346492 387592
rect 346447 387552 346492 387580
rect 346486 387540 346492 387552
rect 346544 387540 346550 387592
rect 346578 387540 346584 387592
rect 346636 387580 346642 387592
rect 354646 387580 354674 387620
rect 450446 387580 450452 387592
rect 346636 387552 346729 387580
rect 354646 387552 450452 387580
rect 346636 387540 346642 387552
rect 450446 387540 450452 387552
rect 450504 387540 450510 387592
rect 346596 387512 346624 387540
rect 407390 387512 407396 387524
rect 346596 387484 407396 387512
rect 407390 387472 407396 387484
rect 407448 387472 407454 387524
rect 346302 387444 346308 387456
rect 346263 387416 346308 387444
rect 346302 387404 346308 387416
rect 346360 387404 346366 387456
rect 412266 387172 412272 387184
rect 373966 387144 412272 387172
rect 367738 387104 367744 387116
rect 367699 387076 367744 387104
rect 367738 387064 367744 387076
rect 367796 387064 367802 387116
rect 367833 387107 367891 387113
rect 367833 387073 367845 387107
rect 367879 387104 367891 387107
rect 371234 387104 371240 387116
rect 367879 387076 371240 387104
rect 367879 387073 367891 387076
rect 367833 387067 367891 387073
rect 371234 387064 371240 387076
rect 371292 387064 371298 387116
rect 22094 386996 22100 387048
rect 22152 387036 22158 387048
rect 367465 387039 367523 387045
rect 367465 387036 367477 387039
rect 22152 387008 367477 387036
rect 22152 386996 22158 387008
rect 367465 387005 367477 387008
rect 367511 387005 367523 387039
rect 367756 387036 367784 387064
rect 368382 387036 368388 387048
rect 367756 387008 368388 387036
rect 367465 386999 367523 387005
rect 368382 386996 368388 387008
rect 368440 387036 368446 387048
rect 373966 387036 373994 387144
rect 412266 387132 412272 387144
rect 412324 387132 412330 387184
rect 368440 387008 373994 387036
rect 368440 386996 368446 387008
rect 367554 386968 367560 386980
rect 367467 386940 367560 386968
rect 367554 386928 367560 386940
rect 367612 386968 367618 386980
rect 367612 386940 373994 386968
rect 367612 386928 367618 386940
rect 368014 386900 368020 386912
rect 367975 386872 368020 386900
rect 368014 386860 368020 386872
rect 368072 386860 368078 386912
rect 373966 386900 373994 386940
rect 450630 386900 450636 386912
rect 373966 386872 450636 386900
rect 450630 386860 450636 386872
rect 450688 386860 450694 386912
rect 353938 384956 353944 385008
rect 353996 384996 354002 385008
rect 495434 384996 495440 385008
rect 353996 384968 495440 384996
rect 353996 384956 354002 384968
rect 495434 384956 495440 384968
rect 495492 384956 495498 385008
rect 95970 384752 95976 384804
rect 96028 384792 96034 384804
rect 199381 384795 199439 384801
rect 199381 384792 199393 384795
rect 96028 384764 199393 384792
rect 96028 384752 96034 384764
rect 199381 384761 199393 384764
rect 199427 384761 199439 384795
rect 199381 384755 199439 384761
rect 108298 384724 108304 384736
rect 108259 384696 108304 384724
rect 108298 384684 108304 384696
rect 108356 384684 108362 384736
rect 89438 384520 89444 384532
rect 89399 384492 89444 384520
rect 89438 384480 89444 384492
rect 89496 384520 89502 384532
rect 89496 384492 93854 384520
rect 89496 384480 89502 384492
rect 93826 384452 93854 384492
rect 414382 384452 414388 384464
rect 93826 384424 414388 384452
rect 414382 384412 414388 384424
rect 414440 384412 414446 384464
rect 89254 384384 89260 384396
rect 89215 384356 89260 384384
rect 89254 384344 89260 384356
rect 89312 384344 89318 384396
rect 142430 384384 142436 384396
rect 103348 384356 142436 384384
rect 103348 384325 103376 384356
rect 142430 384344 142436 384356
rect 142488 384344 142494 384396
rect 103333 384319 103391 384325
rect 103333 384285 103345 384319
rect 103379 384285 103391 384319
rect 103333 384279 103391 384285
rect 103425 384319 103483 384325
rect 103425 384285 103437 384319
rect 103471 384316 103483 384319
rect 132586 384316 132592 384328
rect 103471 384288 122834 384316
rect 132547 384288 132592 384316
rect 103471 384285 103483 384288
rect 103425 384279 103483 384285
rect 88794 384248 88800 384260
rect 88755 384220 88800 384248
rect 88794 384208 88800 384220
rect 88852 384208 88858 384260
rect 122806 384248 122834 384288
rect 132586 384276 132592 384288
rect 132644 384276 132650 384328
rect 403802 384316 403808 384328
rect 142126 384288 403808 384316
rect 142126 384248 142154 384288
rect 403802 384276 403808 384288
rect 403860 384276 403866 384328
rect 122806 384220 142154 384248
rect 200482 384208 200488 384260
rect 200540 384248 200546 384260
rect 232682 384248 232688 384260
rect 200540 384220 232688 384248
rect 200540 384208 200546 384220
rect 232682 384208 232688 384220
rect 232740 384208 232746 384260
rect 89070 384180 89076 384192
rect 89031 384152 89076 384180
rect 89070 384140 89076 384152
rect 89128 384140 89134 384192
rect 89162 384140 89168 384192
rect 89220 384180 89226 384192
rect 89220 384152 89265 384180
rect 89220 384140 89226 384152
rect 103514 384140 103520 384192
rect 103572 384180 103578 384192
rect 132402 384180 132408 384192
rect 103572 384152 103617 384180
rect 132363 384152 132408 384180
rect 103572 384140 103578 384152
rect 132402 384140 132408 384152
rect 132460 384140 132466 384192
rect 198001 384183 198059 384189
rect 198001 384149 198013 384183
rect 198047 384180 198059 384183
rect 200577 384183 200635 384189
rect 200577 384180 200589 384183
rect 198047 384152 200589 384180
rect 198047 384149 198059 384152
rect 198001 384143 198059 384149
rect 200577 384149 200589 384152
rect 200623 384149 200635 384183
rect 200577 384143 200635 384149
rect 177022 383976 177028 383988
rect 176983 383948 177028 383976
rect 177022 383936 177028 383948
rect 177080 383936 177086 383988
rect 259178 383976 259184 383988
rect 177224 383948 259184 383976
rect 177224 383852 177252 383948
rect 259178 383936 259184 383948
rect 259236 383936 259242 383988
rect 198001 383911 198059 383917
rect 198001 383908 198013 383911
rect 177592 383880 198013 383908
rect 177206 383840 177212 383852
rect 177167 383812 177212 383840
rect 177206 383800 177212 383812
rect 177264 383800 177270 383852
rect 177298 383800 177304 383852
rect 177356 383840 177362 383852
rect 177592 383849 177620 383880
rect 198001 383877 198013 383880
rect 198047 383877 198059 383911
rect 198001 383871 198059 383877
rect 200025 383911 200083 383917
rect 200025 383877 200037 383911
rect 200071 383908 200083 383911
rect 200577 383911 200635 383917
rect 200071 383880 200160 383908
rect 200071 383877 200083 383880
rect 200025 383871 200083 383877
rect 177577 383843 177635 383849
rect 177356 383812 177401 383840
rect 177356 383800 177362 383812
rect 177577 383809 177589 383843
rect 177623 383809 177635 383843
rect 199654 383840 199660 383852
rect 177577 383803 177635 383809
rect 180766 383812 199660 383840
rect 177316 383772 177344 383800
rect 180766 383772 180794 383812
rect 199654 383800 199660 383812
rect 199712 383800 199718 383852
rect 199933 383843 199991 383849
rect 199933 383840 199945 383843
rect 199856 383812 199945 383840
rect 177316 383744 180794 383772
rect 199746 383732 199752 383784
rect 199804 383772 199810 383784
rect 199856 383772 199884 383812
rect 199933 383809 199945 383812
rect 199979 383809 199991 383843
rect 200132 383840 200160 383880
rect 200577 383877 200589 383911
rect 200623 383908 200635 383911
rect 279602 383908 279608 383920
rect 200623 383880 279608 383908
rect 200623 383877 200635 383880
rect 200577 383871 200635 383877
rect 279602 383868 279608 383880
rect 279660 383868 279666 383920
rect 200393 383843 200451 383849
rect 200132 383812 200344 383840
rect 199933 383803 199991 383809
rect 199804 383744 199884 383772
rect 199804 383732 199810 383744
rect 200114 383732 200120 383784
rect 200172 383772 200178 383784
rect 200316 383772 200344 383812
rect 200393 383809 200405 383843
rect 200439 383840 200451 383843
rect 334066 383840 334072 383852
rect 200439 383812 334072 383840
rect 200439 383809 200451 383812
rect 200393 383803 200451 383809
rect 334066 383800 334072 383812
rect 334124 383800 334130 383852
rect 311986 383772 311992 383784
rect 200172 383744 200217 383772
rect 200316 383744 311992 383772
rect 200172 383732 200178 383744
rect 311986 383732 311992 383744
rect 312044 383732 312050 383784
rect 177485 383707 177543 383713
rect 177485 383673 177497 383707
rect 177531 383704 177543 383707
rect 317046 383704 317052 383716
rect 177531 383676 317052 383704
rect 177531 383673 177543 383676
rect 177485 383667 177543 383673
rect 317046 383664 317052 383676
rect 317104 383664 317110 383716
rect 199381 383639 199439 383645
rect 199381 383605 199393 383639
rect 199427 383636 199439 383639
rect 199565 383639 199623 383645
rect 199565 383636 199577 383639
rect 199427 383608 199577 383636
rect 199427 383605 199439 383608
rect 199381 383599 199439 383605
rect 199565 383605 199577 383608
rect 199611 383605 199623 383639
rect 199565 383599 199623 383605
rect 199654 383596 199660 383648
rect 199712 383636 199718 383648
rect 200393 383639 200451 383645
rect 200393 383636 200405 383639
rect 199712 383608 200405 383636
rect 199712 383596 199718 383608
rect 200393 383605 200405 383608
rect 200439 383605 200451 383639
rect 200393 383599 200451 383605
rect 13722 383188 13728 383240
rect 13780 383228 13786 383240
rect 96341 383231 96399 383237
rect 96341 383228 96353 383231
rect 13780 383200 96353 383228
rect 13780 383188 13786 383200
rect 96341 383197 96353 383200
rect 96387 383197 96399 383231
rect 130378 383228 130384 383240
rect 130339 383200 130384 383228
rect 96341 383191 96399 383197
rect 130378 383188 130384 383200
rect 130436 383188 130442 383240
rect 322290 383228 322296 383240
rect 322251 383200 322296 383228
rect 322290 383188 322296 383200
rect 322348 383188 322354 383240
rect 136542 381488 136548 381540
rect 136600 381528 136606 381540
rect 464338 381528 464344 381540
rect 136600 381500 464344 381528
rect 136600 381488 136606 381500
rect 464338 381488 464344 381500
rect 464396 381488 464402 381540
rect 39390 381012 39396 381064
rect 39448 381052 39454 381064
rect 40773 381055 40831 381061
rect 39448 381024 40724 381052
rect 39448 381012 39454 381024
rect 40506 380987 40564 380993
rect 40506 380953 40518 380987
rect 40552 380953 40564 380987
rect 40506 380947 40564 380953
rect 39390 380916 39396 380928
rect 39351 380888 39396 380916
rect 39390 380876 39396 380888
rect 39448 380876 39454 380928
rect 40512 380916 40540 380947
rect 40586 380916 40592 380928
rect 40512 380888 40592 380916
rect 40586 380876 40592 380888
rect 40644 380876 40650 380928
rect 40696 380916 40724 381024
rect 40773 381021 40785 381055
rect 40819 381052 40831 381055
rect 89254 381052 89260 381064
rect 40819 381024 89260 381052
rect 40819 381021 40831 381024
rect 40773 381015 40831 381021
rect 89254 381012 89260 381024
rect 89312 381012 89318 381064
rect 136082 380916 136088 380928
rect 40696 380888 136088 380916
rect 136082 380876 136088 380888
rect 136140 380916 136146 380928
rect 136542 380916 136548 380928
rect 136140 380888 136548 380916
rect 136140 380876 136146 380888
rect 136542 380876 136548 380888
rect 136600 380876 136606 380928
rect 274450 380440 274456 380452
rect 274411 380412 274456 380440
rect 274450 380400 274456 380412
rect 274508 380400 274514 380452
rect 70872 378916 74534 378944
rect 70872 378885 70900 378916
rect 70673 378879 70731 378885
rect 70673 378845 70685 378879
rect 70719 378845 70731 378879
rect 70673 378839 70731 378845
rect 70857 378879 70915 378885
rect 70857 378845 70869 378879
rect 70903 378845 70915 378879
rect 71866 378876 71872 378888
rect 71827 378848 71872 378876
rect 70857 378839 70915 378845
rect 70688 378808 70716 378839
rect 71866 378836 71872 378848
rect 71924 378836 71930 378888
rect 74506 378876 74534 378916
rect 259546 378876 259552 378888
rect 74506 378848 259552 378876
rect 259546 378836 259552 378848
rect 259604 378836 259610 378888
rect 71317 378811 71375 378817
rect 71317 378808 71329 378811
rect 70688 378780 71329 378808
rect 71317 378777 71329 378780
rect 71363 378777 71375 378811
rect 71884 378808 71912 378836
rect 95786 378808 95792 378820
rect 71884 378780 95792 378808
rect 71317 378771 71375 378777
rect 95786 378768 95792 378780
rect 95844 378768 95850 378820
rect 70578 378740 70584 378752
rect 70539 378712 70584 378740
rect 70578 378700 70584 378712
rect 70636 378700 70642 378752
rect 309686 375816 309692 375828
rect 309647 375788 309692 375816
rect 309686 375776 309692 375788
rect 309744 375776 309750 375828
rect 308306 375680 308312 375692
rect 308267 375652 308312 375680
rect 308306 375640 308312 375652
rect 308364 375640 308370 375692
rect 5350 375572 5356 375624
rect 5408 375612 5414 375624
rect 207569 375615 207627 375621
rect 207569 375612 207581 375615
rect 5408 375584 207581 375612
rect 5408 375572 5414 375584
rect 207569 375581 207581 375584
rect 207615 375581 207627 375615
rect 308324 375612 308352 375640
rect 342254 375612 342260 375624
rect 308324 375584 342260 375612
rect 207569 375575 207627 375581
rect 342254 375572 342260 375584
rect 342312 375572 342318 375624
rect 8846 375504 8852 375556
rect 8904 375544 8910 375556
rect 308554 375547 308612 375553
rect 308554 375544 308566 375547
rect 8904 375516 308566 375544
rect 8904 375504 8910 375516
rect 308554 375513 308566 375516
rect 308600 375513 308612 375547
rect 308554 375507 308612 375513
rect 309686 375436 309692 375488
rect 309744 375476 309750 375488
rect 366726 375476 366732 375488
rect 309744 375448 366732 375476
rect 309744 375436 309750 375448
rect 366726 375436 366732 375448
rect 366784 375436 366790 375488
rect 409414 375136 409420 375148
rect 409375 375108 409420 375136
rect 409414 375096 409420 375108
rect 409472 375096 409478 375148
rect 404998 375028 405004 375080
rect 405056 375068 405062 375080
rect 409509 375071 409567 375077
rect 409509 375068 409521 375071
rect 405056 375040 409521 375068
rect 405056 375028 405062 375040
rect 409509 375037 409521 375040
rect 409555 375037 409567 375071
rect 409509 375031 409567 375037
rect 409598 375028 409604 375080
rect 409656 375068 409662 375080
rect 419074 375068 419080 375080
rect 409656 375040 419080 375068
rect 409656 375028 409662 375040
rect 419074 375028 419080 375040
rect 419132 375028 419138 375080
rect 409046 374932 409052 374944
rect 409007 374904 409052 374932
rect 409046 374892 409052 374904
rect 409104 374892 409110 374944
rect 95602 374728 95608 374740
rect 95563 374700 95608 374728
rect 95602 374688 95608 374700
rect 95660 374688 95666 374740
rect 450446 374728 450452 374740
rect 450407 374700 450452 374728
rect 450446 374688 450452 374700
rect 450504 374688 450510 374740
rect 95970 374592 95976 374604
rect 95931 374564 95976 374592
rect 95970 374552 95976 374564
rect 96028 374552 96034 374604
rect 95786 374524 95792 374536
rect 95699 374496 95792 374524
rect 95786 374484 95792 374496
rect 95844 374524 95850 374536
rect 152366 374524 152372 374536
rect 95844 374496 152372 374524
rect 95844 374484 95850 374496
rect 152366 374484 152372 374496
rect 152424 374484 152430 374536
rect 450630 374524 450636 374536
rect 450591 374496 450636 374524
rect 450630 374484 450636 374496
rect 450688 374484 450694 374536
rect 441982 372348 441988 372360
rect 441943 372320 441988 372348
rect 441982 372308 441988 372320
rect 442040 372308 442046 372360
rect 233694 371872 233700 371884
rect 233655 371844 233700 371872
rect 233694 371832 233700 371844
rect 233752 371832 233758 371884
rect 233786 371668 233792 371680
rect 233699 371640 233792 371668
rect 233786 371628 233792 371640
rect 233844 371668 233850 371680
rect 366818 371668 366824 371680
rect 233844 371640 366824 371668
rect 233844 371628 233850 371640
rect 366818 371628 366824 371640
rect 366876 371628 366882 371680
rect 214742 370172 214748 370184
rect 214703 370144 214748 370172
rect 214742 370132 214748 370144
rect 214800 370132 214806 370184
rect 335630 369152 335636 369164
rect 325666 369124 335636 369152
rect 293678 369084 293684 369096
rect 293639 369056 293684 369084
rect 293678 369044 293684 369056
rect 293736 369084 293742 369096
rect 325510 369084 325516 369096
rect 293736 369056 325516 369084
rect 293736 369044 293742 369056
rect 325510 369044 325516 369056
rect 325568 369084 325574 369096
rect 325666 369084 325694 369124
rect 335630 369112 335636 369124
rect 335688 369112 335694 369164
rect 325568 369056 325694 369084
rect 325568 369044 325574 369056
rect 293773 368951 293831 368957
rect 293773 368917 293785 368951
rect 293819 368948 293831 368951
rect 311618 368948 311624 368960
rect 293819 368920 311624 368948
rect 293819 368917 293831 368920
rect 293773 368911 293831 368917
rect 311618 368908 311624 368920
rect 311676 368908 311682 368960
rect 2774 366664 2780 366716
rect 2832 366704 2838 366716
rect 4706 366704 4712 366716
rect 2832 366676 4712 366704
rect 2832 366664 2838 366676
rect 4706 366664 4712 366676
rect 4764 366664 4770 366716
rect 360562 366568 360568 366580
rect 360523 366540 360568 366568
rect 360562 366528 360568 366540
rect 360620 366528 360626 366580
rect 360378 366432 360384 366444
rect 360339 366404 360384 366432
rect 360378 366392 360384 366404
rect 360436 366392 360442 366444
rect 360194 366364 360200 366376
rect 360155 366336 360200 366364
rect 360194 366324 360200 366336
rect 360252 366324 360258 366376
rect 314562 365712 314568 365764
rect 314620 365752 314626 365764
rect 495434 365752 495440 365764
rect 314620 365724 495440 365752
rect 314620 365712 314626 365724
rect 495434 365712 495440 365724
rect 495492 365712 495498 365764
rect 143445 365483 143503 365489
rect 143445 365449 143457 365483
rect 143491 365480 143503 365483
rect 473722 365480 473728 365492
rect 143491 365452 151814 365480
rect 473683 365452 473728 365480
rect 143491 365449 143503 365452
rect 143445 365443 143503 365449
rect 142985 365415 143043 365421
rect 142985 365381 142997 365415
rect 143031 365412 143043 365415
rect 143074 365412 143080 365424
rect 143031 365384 143080 365412
rect 143031 365381 143043 365384
rect 142985 365375 143043 365381
rect 143074 365372 143080 365384
rect 143132 365372 143138 365424
rect 143169 365415 143227 365421
rect 143169 365381 143181 365415
rect 143215 365412 143227 365415
rect 151786 365412 151814 365452
rect 473722 365440 473728 365452
rect 473780 365440 473786 365492
rect 263870 365412 263876 365424
rect 143215 365384 149560 365412
rect 151786 365384 263876 365412
rect 143215 365381 143227 365384
rect 143169 365375 143227 365381
rect 143353 365347 143411 365353
rect 143353 365313 143365 365347
rect 143399 365344 143411 365347
rect 143445 365347 143503 365353
rect 143445 365344 143457 365347
rect 143399 365316 143457 365344
rect 143399 365313 143411 365316
rect 143353 365307 143411 365313
rect 143445 365313 143457 365316
rect 143491 365313 143503 365347
rect 149532 365344 149560 365384
rect 263870 365372 263876 365384
rect 263928 365372 263934 365424
rect 264054 365344 264060 365356
rect 149532 365316 264060 365344
rect 143445 365307 143503 365313
rect 264054 365304 264060 365316
rect 264112 365304 264118 365356
rect 473630 365344 473636 365356
rect 473591 365316 473636 365344
rect 473630 365304 473636 365316
rect 473688 365304 473694 365356
rect 143074 365100 143080 365152
rect 143132 365140 143138 365152
rect 355594 365140 355600 365152
rect 143132 365112 355600 365140
rect 143132 365100 143138 365112
rect 355594 365100 355600 365112
rect 355652 365100 355658 365152
rect 470410 364732 470416 364744
rect 470323 364704 470416 364732
rect 470410 364692 470416 364704
rect 470468 364732 470474 364744
rect 486970 364732 486976 364744
rect 470468 364704 486976 364732
rect 470468 364692 470474 364704
rect 486970 364692 486976 364704
rect 487028 364692 487034 364744
rect 248138 364624 248144 364676
rect 248196 364664 248202 364676
rect 470658 364667 470716 364673
rect 470658 364664 470670 364667
rect 248196 364636 470670 364664
rect 248196 364624 248202 364636
rect 470658 364633 470670 364636
rect 470704 364633 470716 364667
rect 470658 364627 470716 364633
rect 471793 364599 471851 364605
rect 471793 364565 471805 364599
rect 471839 364596 471851 364599
rect 496354 364596 496360 364608
rect 471839 364568 496360 364596
rect 471839 364565 471851 364568
rect 471793 364559 471851 364565
rect 496354 364556 496360 364568
rect 496412 364556 496418 364608
rect 153010 362584 153016 362636
rect 153068 362624 153074 362636
rect 180426 362624 180432 362636
rect 153068 362596 180288 362624
rect 180387 362596 180432 362624
rect 153068 362584 153074 362596
rect 180260 362565 180288 362596
rect 180426 362584 180432 362596
rect 180484 362584 180490 362636
rect 49881 362559 49939 362565
rect 49881 362525 49893 362559
rect 49927 362556 49939 362559
rect 180245 362559 180303 362565
rect 49927 362528 161474 362556
rect 49927 362525 49939 362528
rect 49881 362519 49939 362525
rect 161446 362420 161474 362528
rect 180245 362525 180257 362559
rect 180291 362525 180303 362559
rect 316034 362556 316040 362568
rect 180245 362519 180303 362525
rect 180766 362528 316040 362556
rect 180058 362488 180064 362500
rect 180019 362460 180064 362488
rect 180058 362448 180064 362460
rect 180116 362448 180122 362500
rect 180766 362420 180794 362528
rect 316034 362516 316040 362528
rect 316092 362516 316098 362568
rect 161446 362392 180794 362420
rect 426986 361564 426992 361616
rect 427044 361604 427050 361616
rect 495434 361604 495440 361616
rect 427044 361576 495440 361604
rect 427044 361564 427050 361576
rect 495434 361564 495440 361576
rect 495492 361564 495498 361616
rect 244366 360380 244372 360392
rect 244327 360352 244372 360380
rect 244366 360340 244372 360352
rect 244424 360340 244430 360392
rect 402790 360380 402796 360392
rect 402751 360352 402796 360380
rect 402790 360340 402796 360352
rect 402848 360340 402854 360392
rect 402974 360340 402980 360392
rect 403032 360380 403038 360392
rect 403032 360352 403077 360380
rect 403032 360340 403038 360352
rect 336182 360204 336188 360256
rect 336240 360244 336246 360256
rect 402885 360247 402943 360253
rect 402885 360244 402897 360247
rect 336240 360216 402897 360244
rect 336240 360204 336246 360216
rect 402885 360213 402897 360216
rect 402931 360213 402943 360247
rect 402885 360207 402943 360213
rect 361482 359904 361488 359916
rect 361443 359876 361488 359904
rect 361482 359864 361488 359876
rect 361540 359904 361546 359916
rect 468018 359904 468024 359916
rect 361540 359876 468024 359904
rect 361540 359864 361546 359876
rect 468018 359864 468024 359876
rect 468076 359864 468082 359916
rect 361666 359700 361672 359712
rect 361627 359672 361672 359700
rect 361666 359660 361672 359672
rect 361724 359700 361730 359712
rect 434898 359700 434904 359712
rect 361724 359672 434904 359700
rect 361724 359660 361730 359672
rect 434898 359660 434904 359672
rect 434956 359660 434962 359712
rect 88334 359360 88340 359372
rect 88295 359332 88340 359360
rect 88334 359320 88340 359332
rect 88392 359320 88398 359372
rect 88153 359295 88211 359301
rect 88153 359261 88165 359295
rect 88199 359292 88211 359295
rect 93486 359292 93492 359304
rect 88199 359264 93492 359292
rect 88199 359261 88211 359264
rect 88153 359255 88211 359261
rect 93486 359252 93492 359264
rect 93544 359252 93550 359304
rect 87969 359159 88027 359165
rect 87969 359125 87981 359159
rect 88015 359156 88027 359159
rect 312538 359156 312544 359168
rect 88015 359128 312544 359156
rect 88015 359125 88027 359128
rect 87969 359119 88027 359125
rect 312538 359116 312544 359128
rect 312596 359116 312602 359168
rect 90634 356776 90640 356788
rect 90595 356748 90640 356776
rect 90634 356736 90640 356748
rect 90692 356736 90698 356788
rect 89254 356668 89260 356720
rect 89312 356708 89318 356720
rect 89312 356680 93854 356708
rect 89312 356668 89318 356680
rect 56686 356600 56692 356652
rect 56744 356640 56750 356652
rect 89513 356643 89571 356649
rect 89513 356640 89525 356643
rect 56744 356612 89525 356640
rect 56744 356600 56750 356612
rect 89513 356609 89525 356612
rect 89559 356609 89571 356643
rect 93826 356640 93854 356680
rect 106366 356640 106372 356652
rect 93826 356612 106372 356640
rect 89513 356603 89571 356609
rect 106366 356600 106372 356612
rect 106424 356600 106430 356652
rect 89254 356572 89260 356584
rect 89215 356544 89260 356572
rect 89254 356532 89260 356544
rect 89312 356532 89318 356584
rect 3786 356056 3792 356108
rect 3844 356096 3850 356108
rect 200025 356099 200083 356105
rect 200025 356096 200037 356099
rect 3844 356068 200037 356096
rect 3844 356056 3850 356068
rect 200025 356065 200037 356068
rect 200071 356065 200083 356099
rect 200025 356059 200083 356065
rect 7469 356031 7527 356037
rect 7469 355997 7481 356031
rect 7515 356028 7527 356031
rect 67082 356028 67088 356040
rect 7515 356000 67088 356028
rect 7515 355997 7527 356000
rect 7469 355991 7527 355997
rect 67082 355988 67088 356000
rect 67140 355988 67146 356040
rect 361574 356028 361580 356040
rect 361487 356000 361580 356028
rect 361574 355988 361580 356000
rect 361632 356028 361638 356040
rect 402422 356028 402428 356040
rect 361632 356000 402428 356028
rect 361632 355988 361638 356000
rect 402422 355988 402428 356000
rect 402480 355988 402486 356040
rect 7377 355895 7435 355901
rect 7377 355861 7389 355895
rect 7423 355892 7435 355895
rect 67542 355892 67548 355904
rect 7423 355864 67548 355892
rect 7423 355861 7435 355864
rect 7377 355855 7435 355861
rect 67542 355852 67548 355864
rect 67600 355852 67606 355904
rect 220538 355852 220544 355904
rect 220596 355892 220602 355904
rect 361393 355895 361451 355901
rect 361393 355892 361405 355895
rect 220596 355864 361405 355892
rect 220596 355852 220602 355864
rect 361393 355861 361405 355864
rect 361439 355861 361451 355895
rect 361393 355855 361451 355861
rect 67542 355308 67548 355360
rect 67600 355348 67606 355360
rect 207014 355348 207020 355360
rect 67600 355320 207020 355348
rect 67600 355308 67606 355320
rect 207014 355308 207020 355320
rect 207072 355308 207078 355360
rect 326982 355308 326988 355360
rect 327040 355348 327046 355360
rect 403713 355351 403771 355357
rect 403713 355348 403725 355351
rect 327040 355320 403725 355348
rect 327040 355308 327046 355320
rect 403713 355317 403725 355320
rect 403759 355317 403771 355351
rect 403713 355311 403771 355317
rect 195057 354399 195115 354405
rect 195057 354365 195069 354399
rect 195103 354396 195115 354399
rect 195238 354396 195244 354408
rect 195103 354368 195244 354396
rect 195103 354365 195115 354368
rect 195057 354359 195115 354365
rect 195238 354356 195244 354368
rect 195296 354396 195302 354408
rect 195422 354396 195428 354408
rect 195296 354368 195428 354396
rect 195296 354356 195302 354368
rect 195422 354356 195428 354368
rect 195480 354356 195486 354408
rect 193674 354220 193680 354272
rect 193732 354260 193738 354272
rect 194413 354263 194471 354269
rect 194413 354260 194425 354263
rect 193732 354232 194425 354260
rect 193732 354220 193738 354232
rect 194413 354229 194425 354232
rect 194459 354229 194471 354263
rect 194413 354223 194471 354229
rect 194137 353855 194195 353861
rect 194137 353821 194149 353855
rect 194183 353852 194195 353855
rect 195885 353855 195943 353861
rect 195885 353852 195897 353855
rect 194183 353824 195897 353852
rect 194183 353821 194195 353824
rect 194137 353815 194195 353821
rect 195885 353821 195897 353824
rect 195931 353852 195943 353855
rect 296070 353852 296076 353864
rect 195931 353824 296076 353852
rect 195931 353821 195943 353824
rect 195885 353815 195943 353821
rect 296070 353812 296076 353824
rect 296128 353812 296134 353864
rect 54018 353744 54024 353796
rect 54076 353784 54082 353796
rect 194781 353787 194839 353793
rect 194781 353784 194793 353787
rect 54076 353756 194793 353784
rect 54076 353744 54082 353756
rect 194781 353753 194793 353756
rect 194827 353753 194839 353787
rect 194781 353747 194839 353753
rect 193677 353719 193735 353725
rect 193677 353685 193689 353719
rect 193723 353716 193735 353719
rect 193723 353688 194272 353716
rect 193723 353685 193735 353688
rect 193677 353679 193735 353685
rect 193582 353376 193588 353388
rect 193543 353348 193588 353376
rect 193582 353336 193588 353348
rect 193640 353336 193646 353388
rect 193674 353336 193680 353388
rect 193732 353376 193738 353388
rect 193953 353379 194011 353385
rect 193732 353348 193777 353376
rect 193732 353336 193738 353348
rect 193953 353345 193965 353379
rect 193999 353376 194011 353379
rect 194244 353376 194272 353688
rect 194594 353444 194600 353456
rect 194555 353416 194600 353444
rect 194594 353404 194600 353416
rect 194652 353404 194658 353456
rect 195422 353376 195428 353388
rect 193999 353348 194272 353376
rect 195335 353348 195428 353376
rect 193999 353345 194011 353348
rect 193953 353339 194011 353345
rect 195422 353336 195428 353348
rect 195480 353376 195486 353388
rect 323578 353376 323584 353388
rect 195480 353348 323584 353376
rect 195480 353336 195486 353348
rect 323578 353336 323584 353348
rect 323636 353336 323642 353388
rect 106182 353268 106188 353320
rect 106240 353308 106246 353320
rect 193401 353311 193459 353317
rect 193401 353308 193413 353311
rect 106240 353280 193413 353308
rect 106240 353268 106246 353280
rect 193401 353277 193413 353280
rect 193447 353277 193459 353311
rect 193858 353308 193864 353320
rect 193819 353280 193864 353308
rect 193401 353271 193459 353277
rect 193858 353268 193864 353280
rect 193916 353268 193922 353320
rect 141053 351679 141111 351685
rect 141053 351645 141065 351679
rect 141099 351676 141111 351679
rect 366358 351676 366364 351688
rect 141099 351648 366364 351676
rect 141099 351645 141111 351648
rect 141053 351639 141111 351645
rect 366358 351636 366364 351648
rect 366416 351636 366422 351688
rect 451458 349500 451464 349512
rect 451419 349472 451464 349500
rect 451458 349460 451464 349472
rect 451516 349460 451522 349512
rect 9398 349324 9404 349376
rect 9456 349364 9462 349376
rect 451553 349367 451611 349373
rect 451553 349364 451565 349367
rect 9456 349336 451565 349364
rect 9456 349324 9462 349336
rect 451553 349333 451565 349336
rect 451599 349333 451611 349367
rect 451553 349327 451611 349333
rect 99834 349052 99840 349104
rect 99892 349092 99898 349104
rect 100662 349092 100668 349104
rect 99892 349064 100668 349092
rect 99892 349052 99898 349064
rect 100662 349052 100668 349064
rect 100720 349052 100726 349104
rect 5353 348619 5411 348625
rect 5353 348616 5365 348619
rect 4816 348588 5365 348616
rect 4709 348415 4767 348421
rect 4709 348381 4721 348415
rect 4755 348412 4767 348415
rect 4816 348412 4844 348588
rect 5353 348585 5365 348588
rect 5399 348585 5411 348619
rect 5353 348579 5411 348585
rect 99834 348548 99840 348560
rect 4908 348520 99840 348548
rect 4908 348421 4936 348520
rect 99834 348508 99840 348520
rect 99892 348508 99898 348560
rect 5353 348483 5411 348489
rect 5353 348449 5365 348483
rect 5399 348480 5411 348483
rect 99650 348480 99656 348492
rect 5399 348452 99656 348480
rect 5399 348449 5411 348452
rect 5353 348443 5411 348449
rect 99650 348440 99656 348452
rect 99708 348440 99714 348492
rect 5092 348421 5212 348422
rect 4755 348384 4844 348412
rect 4893 348415 4951 348421
rect 4755 348381 4767 348384
rect 4709 348375 4767 348381
rect 4893 348381 4905 348415
rect 4939 348381 4951 348415
rect 4893 348375 4951 348381
rect 4985 348415 5043 348421
rect 4985 348381 4997 348415
rect 5031 348381 5043 348415
rect 4985 348375 5043 348381
rect 5078 348415 5212 348421
rect 5078 348381 5090 348415
rect 5124 348394 5212 348415
rect 5124 348381 5136 348394
rect 5078 348375 5136 348381
rect 4614 348276 4620 348288
rect 4575 348248 4620 348276
rect 4614 348236 4620 348248
rect 4672 348236 4678 348288
rect 5000 348276 5028 348375
rect 5184 348344 5212 348394
rect 5261 348415 5319 348421
rect 5261 348381 5273 348415
rect 5307 348412 5319 348415
rect 470594 348412 470600 348424
rect 5307 348384 470600 348412
rect 5307 348381 5319 348384
rect 5261 348375 5319 348381
rect 470594 348372 470600 348384
rect 470652 348372 470658 348424
rect 232314 348344 232320 348356
rect 5184 348316 232320 348344
rect 232314 348304 232320 348316
rect 232372 348304 232378 348356
rect 100938 348276 100944 348288
rect 5000 348248 100944 348276
rect 100938 348236 100944 348248
rect 100996 348236 101002 348288
rect 485406 346848 485412 346860
rect 485367 346820 485412 346848
rect 485406 346808 485412 346820
rect 485464 346808 485470 346860
rect 485590 346848 485596 346860
rect 485551 346820 485596 346848
rect 485590 346808 485596 346820
rect 485648 346808 485654 346860
rect 420914 346604 420920 346656
rect 420972 346644 420978 346656
rect 485501 346647 485559 346653
rect 485501 346644 485513 346647
rect 420972 346616 485513 346644
rect 420972 346604 420978 346616
rect 485501 346613 485513 346616
rect 485547 346613 485559 346647
rect 485501 346607 485559 346613
rect 5258 344428 5264 344480
rect 5316 344468 5322 344480
rect 376205 344471 376263 344477
rect 376205 344468 376217 344471
rect 5316 344440 376217 344468
rect 5316 344428 5322 344440
rect 376205 344437 376217 344440
rect 376251 344437 376263 344471
rect 376205 344431 376263 344437
rect 233326 344264 233332 344276
rect 233287 344236 233332 344264
rect 233326 344224 233332 344236
rect 233384 344224 233390 344276
rect 232682 344128 232688 344140
rect 232643 344100 232688 344128
rect 232682 344088 232688 344100
rect 232740 344128 232746 344140
rect 257062 344128 257068 344140
rect 232740 344100 257068 344128
rect 232740 344088 232746 344100
rect 257062 344088 257068 344100
rect 257120 344088 257126 344140
rect 29549 344063 29607 344069
rect 29549 344029 29561 344063
rect 29595 344060 29607 344063
rect 432598 344060 432604 344072
rect 29595 344032 432604 344060
rect 29595 344029 29607 344032
rect 29549 344023 29607 344029
rect 432598 344020 432604 344032
rect 432656 344020 432662 344072
rect 7926 343884 7932 343936
rect 7984 343924 7990 343936
rect 232869 343927 232927 343933
rect 232869 343924 232881 343927
rect 7984 343896 232881 343924
rect 7984 343884 7990 343896
rect 232869 343893 232881 343896
rect 232915 343893 232927 343927
rect 232869 343887 232927 343893
rect 232958 343884 232964 343936
rect 233016 343924 233022 343936
rect 233016 343896 233061 343924
rect 233016 343884 233022 343896
rect 393222 339668 393228 339720
rect 393280 339708 393286 339720
rect 410981 339711 411039 339717
rect 410981 339708 410993 339711
rect 393280 339680 410993 339708
rect 393280 339668 393286 339680
rect 410981 339677 410993 339680
rect 411027 339677 411039 339711
rect 410981 339671 411039 339677
rect 344738 339232 344744 339244
rect 344651 339204 344744 339232
rect 344738 339192 344744 339204
rect 344796 339232 344802 339244
rect 360378 339232 360384 339244
rect 344796 339204 360384 339232
rect 344796 339192 344802 339204
rect 360378 339192 360384 339204
rect 360436 339192 360442 339244
rect 79778 339124 79784 339176
rect 79836 339164 79842 339176
rect 344557 339167 344615 339173
rect 344557 339164 344569 339167
rect 79836 339136 344569 339164
rect 79836 339124 79842 339136
rect 344557 339133 344569 339136
rect 344603 339133 344615 339167
rect 344557 339127 344615 339133
rect 344922 339028 344928 339040
rect 344883 339000 344928 339028
rect 344922 338988 344928 339000
rect 344980 338988 344986 339040
rect 385126 338144 385132 338156
rect 385087 338116 385132 338144
rect 385126 338104 385132 338116
rect 385184 338104 385190 338156
rect 385218 338104 385224 338156
rect 385276 338144 385282 338156
rect 385276 338116 385321 338144
rect 385276 338104 385282 338116
rect 218977 337739 219035 337745
rect 218977 337705 218989 337739
rect 219023 337736 219035 337739
rect 312262 337736 312268 337748
rect 219023 337708 312268 337736
rect 219023 337705 219035 337708
rect 218977 337699 219035 337705
rect 312262 337696 312268 337708
rect 312320 337696 312326 337748
rect 218793 337603 218851 337609
rect 218793 337600 218805 337603
rect 200086 337572 218805 337600
rect 2958 337492 2964 337544
rect 3016 337532 3022 337544
rect 200086 337532 200114 337572
rect 218793 337569 218805 337572
rect 218839 337600 218851 337603
rect 218839 337572 219434 337600
rect 218839 337569 218851 337572
rect 218793 337563 218851 337569
rect 218698 337532 218704 337544
rect 3016 337504 200114 337532
rect 218659 337504 218704 337532
rect 3016 337492 3022 337504
rect 218698 337492 218704 337504
rect 218756 337492 218762 337544
rect 219406 337532 219434 337572
rect 312354 337532 312360 337544
rect 219406 337504 312360 337532
rect 312354 337492 312360 337504
rect 312412 337532 312418 337544
rect 318794 337532 318800 337544
rect 312412 337504 318800 337532
rect 312412 337492 312418 337504
rect 318794 337492 318800 337504
rect 318852 337492 318858 337544
rect 218977 337467 219035 337473
rect 218977 337433 218989 337467
rect 219023 337464 219035 337467
rect 231026 337464 231032 337476
rect 219023 337436 231032 337464
rect 219023 337433 219035 337436
rect 218977 337427 219035 337433
rect 231026 337424 231032 337436
rect 231084 337464 231090 337476
rect 426894 337464 426900 337476
rect 231084 337436 426900 337464
rect 231084 337424 231090 337436
rect 426894 337424 426900 337436
rect 426952 337424 426958 337476
rect 218514 337396 218520 337408
rect 218475 337368 218520 337396
rect 218514 337356 218520 337368
rect 218572 337396 218578 337408
rect 268746 337396 268752 337408
rect 218572 337368 268752 337396
rect 218572 337356 218578 337368
rect 268746 337356 268752 337368
rect 268804 337356 268810 337408
rect 3142 336676 3148 336728
rect 3200 336716 3206 336728
rect 5350 336716 5356 336728
rect 3200 336688 5356 336716
rect 3200 336676 3206 336688
rect 5350 336676 5356 336688
rect 5408 336676 5414 336728
rect 106182 336104 106188 336116
rect 106108 336076 106188 336104
rect 106108 336045 106136 336076
rect 106182 336064 106188 336076
rect 106240 336064 106246 336116
rect 106102 336039 106160 336045
rect 106102 336005 106114 336039
rect 106148 336005 106160 336039
rect 106102 335999 106160 336005
rect 106366 335968 106372 335980
rect 106327 335940 106372 335968
rect 106366 335928 106372 335940
rect 106424 335968 106430 335980
rect 106424 335940 113174 335968
rect 106424 335928 106430 335940
rect 113146 335900 113174 335940
rect 137922 335900 137928 335912
rect 113146 335872 137928 335900
rect 137922 335860 137928 335872
rect 137980 335860 137986 335912
rect 4062 335724 4068 335776
rect 4120 335764 4126 335776
rect 104989 335767 105047 335773
rect 104989 335764 105001 335767
rect 4120 335736 105001 335764
rect 4120 335724 4126 335736
rect 104989 335733 105001 335736
rect 105035 335764 105047 335767
rect 193582 335764 193588 335776
rect 105035 335736 193588 335764
rect 105035 335733 105047 335736
rect 104989 335727 105047 335733
rect 193582 335724 193588 335736
rect 193640 335724 193646 335776
rect 68189 335359 68247 335365
rect 68189 335325 68201 335359
rect 68235 335356 68247 335359
rect 115934 335356 115940 335368
rect 68235 335328 115940 335356
rect 68235 335325 68247 335328
rect 68189 335319 68247 335325
rect 115934 335316 115940 335328
rect 115992 335316 115998 335368
rect 365806 334676 365812 334688
rect 365767 334648 365812 334676
rect 365806 334636 365812 334648
rect 365864 334636 365870 334688
rect 310606 334364 310612 334416
rect 310664 334404 310670 334416
rect 310664 334376 311894 334404
rect 310664 334364 310670 334376
rect 310885 334339 310943 334345
rect 310885 334305 310897 334339
rect 310931 334336 310943 334339
rect 311713 334339 311771 334345
rect 311713 334336 311725 334339
rect 310931 334308 311725 334336
rect 310931 334305 310943 334308
rect 310885 334299 310943 334305
rect 311713 334305 311725 334308
rect 311759 334305 311771 334339
rect 311866 334336 311894 334376
rect 385218 334336 385224 334348
rect 311866 334308 385224 334336
rect 311713 334299 311771 334305
rect 385218 334296 385224 334308
rect 385276 334296 385282 334348
rect 310606 334268 310612 334280
rect 310567 334240 310612 334268
rect 310606 334228 310612 334240
rect 310664 334228 310670 334280
rect 310790 334268 310796 334280
rect 310751 334240 310796 334268
rect 310790 334228 310796 334240
rect 310848 334228 310854 334280
rect 310978 334268 311036 334274
rect 310978 334234 310990 334268
rect 311024 334234 311036 334268
rect 310978 334228 311036 334234
rect 311161 334271 311219 334277
rect 311161 334237 311173 334271
rect 311207 334268 311219 334271
rect 314657 334271 314715 334277
rect 314657 334268 314669 334271
rect 311207 334240 314669 334268
rect 311207 334237 311219 334240
rect 311161 334231 311219 334237
rect 314657 334237 314669 334240
rect 314703 334237 314715 334271
rect 314657 334231 314715 334237
rect 314749 334271 314807 334277
rect 314749 334237 314761 334271
rect 314795 334268 314807 334271
rect 390922 334268 390928 334280
rect 314795 334240 390928 334268
rect 314795 334237 314807 334240
rect 314749 334231 314807 334237
rect 390922 334228 390928 334240
rect 390980 334228 390986 334280
rect 310993 334200 311021 334228
rect 311066 334200 311072 334212
rect 310979 334172 311072 334200
rect 311066 334160 311072 334172
rect 311124 334200 311130 334212
rect 314473 334203 314531 334209
rect 314473 334200 314485 334203
rect 311124 334172 314485 334200
rect 311124 334160 311130 334172
rect 314473 334169 314485 334172
rect 314519 334169 314531 334203
rect 331766 334200 331772 334212
rect 314473 334163 314531 334169
rect 325666 334172 331772 334200
rect 89070 334092 89076 334144
rect 89128 334132 89134 334144
rect 310517 334135 310575 334141
rect 310517 334132 310529 334135
rect 89128 334104 310529 334132
rect 89128 334092 89134 334104
rect 310517 334101 310529 334104
rect 310563 334101 310575 334135
rect 310517 334095 310575 334101
rect 314657 334067 314715 334073
rect 314657 334033 314669 334067
rect 314703 334064 314715 334067
rect 318150 334064 318156 334076
rect 314703 334036 318156 334064
rect 314703 334033 314715 334036
rect 314657 334027 314715 334033
rect 318150 334024 318156 334036
rect 318208 334024 318214 334076
rect 325666 334064 325694 334172
rect 331766 334160 331772 334172
rect 331824 334160 331830 334212
rect 321526 334036 325694 334064
rect 311713 333999 311771 334005
rect 311713 333965 311725 333999
rect 311759 333996 311771 333999
rect 321526 333996 321554 334036
rect 311759 333968 321554 333996
rect 311759 333965 311771 333968
rect 311713 333959 311771 333965
rect 38838 333248 38844 333260
rect 9600 333220 38844 333248
rect 9600 333189 9628 333220
rect 38838 333208 38844 333220
rect 38896 333208 38902 333260
rect 9585 333183 9643 333189
rect 9585 333149 9597 333183
rect 9631 333149 9643 333183
rect 9585 333143 9643 333149
rect 9861 333183 9919 333189
rect 9861 333149 9873 333183
rect 9907 333180 9919 333183
rect 175550 333180 175556 333192
rect 9907 333152 175556 333180
rect 9907 333149 9919 333152
rect 9861 333143 9919 333149
rect 175550 333140 175556 333152
rect 175608 333140 175614 333192
rect 9309 333115 9367 333121
rect 9309 333081 9321 333115
rect 9355 333112 9367 333115
rect 176010 333112 176016 333124
rect 9355 333084 176016 333112
rect 9355 333081 9367 333084
rect 9309 333075 9367 333081
rect 176010 333072 176016 333084
rect 176068 333072 176074 333124
rect 9122 333004 9128 333056
rect 9180 333044 9186 333056
rect 9493 333047 9551 333053
rect 9493 333044 9505 333047
rect 9180 333016 9505 333044
rect 9180 333004 9186 333016
rect 9493 333013 9505 333016
rect 9539 333013 9551 333047
rect 9493 333007 9551 333013
rect 9677 333047 9735 333053
rect 9677 333013 9689 333047
rect 9723 333044 9735 333047
rect 401134 333044 401140 333056
rect 9723 333016 401140 333044
rect 9723 333013 9735 333016
rect 9677 333007 9735 333013
rect 401134 333004 401140 333016
rect 401192 333004 401198 333056
rect 9122 332800 9128 332852
rect 9180 332840 9186 332852
rect 175734 332840 175740 332852
rect 9180 332812 175740 332840
rect 9180 332800 9186 332812
rect 175734 332800 175740 332812
rect 175792 332800 175798 332852
rect 62209 332639 62267 332645
rect 62209 332605 62221 332639
rect 62255 332636 62267 332639
rect 463694 332636 463700 332648
rect 62255 332608 463700 332636
rect 62255 332605 62267 332608
rect 62209 332599 62267 332605
rect 463694 332596 463700 332608
rect 463752 332596 463758 332648
rect 3602 332528 3608 332580
rect 3660 332568 3666 332580
rect 441982 332568 441988 332580
rect 3660 332540 441988 332568
rect 3660 332528 3666 332540
rect 441982 332528 441988 332540
rect 442040 332528 442046 332580
rect 87785 331415 87843 331421
rect 87785 331381 87797 331415
rect 87831 331412 87843 331415
rect 311250 331412 311256 331424
rect 87831 331384 311256 331412
rect 87831 331381 87843 331384
rect 87785 331375 87843 331381
rect 311250 331372 311256 331384
rect 311308 331372 311314 331424
rect 363506 331208 363512 331220
rect 363467 331180 363512 331208
rect 363506 331168 363512 331180
rect 363564 331168 363570 331220
rect 417510 329780 417516 329792
rect 383626 329752 417516 329780
rect 381541 329579 381599 329585
rect 381541 329545 381553 329579
rect 381587 329545 381599 329579
rect 381541 329539 381599 329545
rect 381633 329579 381691 329585
rect 381633 329545 381645 329579
rect 381679 329576 381691 329579
rect 383626 329576 383654 329752
rect 417510 329740 417516 329752
rect 417568 329780 417574 329792
rect 417786 329780 417792 329792
rect 417568 329752 417792 329780
rect 417568 329740 417574 329752
rect 417786 329740 417792 329752
rect 417844 329740 417850 329792
rect 417878 329576 417884 329588
rect 381679 329548 383654 329576
rect 393286 329548 417884 329576
rect 381679 329545 381691 329548
rect 381633 329539 381691 329545
rect 381556 329508 381584 329539
rect 393286 329508 393314 329548
rect 417878 329536 417884 329548
rect 417936 329536 417942 329588
rect 381556 329480 393314 329508
rect 381446 329440 381452 329452
rect 381407 329412 381452 329440
rect 381446 329400 381452 329412
rect 381504 329400 381510 329452
rect 381817 329443 381875 329449
rect 381817 329409 381829 329443
rect 381863 329440 381875 329443
rect 438302 329440 438308 329452
rect 381863 329412 383654 329440
rect 438263 329412 438308 329440
rect 381863 329409 381875 329412
rect 381817 329403 381875 329409
rect 251177 329375 251235 329381
rect 251177 329341 251189 329375
rect 251223 329372 251235 329375
rect 252373 329375 252431 329381
rect 252373 329372 252385 329375
rect 251223 329344 252385 329372
rect 251223 329341 251235 329344
rect 251177 329335 251235 329341
rect 252373 329341 252385 329344
rect 252419 329341 252431 329375
rect 383626 329372 383654 329412
rect 438302 329400 438308 329412
rect 438360 329400 438366 329452
rect 438486 329440 438492 329452
rect 438447 329412 438492 329440
rect 438486 329400 438492 329412
rect 438544 329400 438550 329452
rect 439958 329372 439964 329384
rect 383626 329344 439964 329372
rect 252373 329335 252431 329341
rect 439958 329332 439964 329344
rect 440016 329332 440022 329384
rect 48222 329264 48228 329316
rect 48280 329304 48286 329316
rect 381265 329307 381323 329313
rect 381265 329304 381277 329307
rect 48280 329276 381277 329304
rect 48280 329264 48286 329276
rect 381265 329273 381277 329276
rect 381311 329273 381323 329307
rect 381265 329267 381323 329273
rect 417510 329264 417516 329316
rect 417568 329304 417574 329316
rect 477678 329304 477684 329316
rect 417568 329276 477684 329304
rect 417568 329264 417574 329276
rect 477678 329264 477684 329276
rect 477736 329264 477742 329316
rect 46198 329196 46204 329248
rect 46256 329236 46262 329248
rect 438397 329239 438455 329245
rect 438397 329236 438409 329239
rect 46256 329208 438409 329236
rect 46256 329196 46262 329208
rect 438397 329205 438409 329208
rect 438443 329205 438455 329239
rect 438397 329199 438455 329205
rect 5258 328992 5264 329044
rect 5316 329032 5322 329044
rect 251177 329035 251235 329041
rect 251177 329032 251189 329035
rect 5316 329004 251189 329032
rect 5316 328992 5322 329004
rect 251177 329001 251189 329004
rect 251223 329001 251235 329035
rect 251177 328995 251235 329001
rect 381446 328992 381452 329044
rect 381504 329032 381510 329044
rect 481726 329032 481732 329044
rect 381504 329004 481732 329032
rect 381504 328992 381510 329004
rect 481726 328992 481732 329004
rect 481784 328992 481790 329044
rect 5166 327700 5172 327752
rect 5224 327740 5230 327752
rect 208489 327743 208547 327749
rect 208489 327740 208501 327743
rect 5224 327712 208501 327740
rect 5224 327700 5230 327712
rect 208489 327709 208501 327712
rect 208535 327709 208547 327743
rect 208489 327703 208547 327709
rect 423766 327360 423772 327412
rect 423824 327400 423830 327412
rect 424045 327403 424103 327409
rect 424045 327400 424057 327403
rect 423824 327372 424057 327400
rect 423824 327360 423830 327372
rect 424045 327369 424057 327372
rect 424091 327369 424103 327403
rect 424045 327363 424103 327369
rect 423950 327264 423956 327276
rect 423911 327236 423956 327264
rect 423950 327224 423956 327236
rect 424008 327224 424014 327276
rect 14458 326612 14464 326664
rect 14516 326652 14522 326664
rect 87049 326655 87107 326661
rect 87049 326652 87061 326655
rect 14516 326624 87061 326652
rect 14516 326612 14522 326624
rect 87049 326621 87061 326624
rect 87095 326621 87107 326655
rect 87049 326615 87107 326621
rect 93302 326176 93308 326188
rect 93263 326148 93308 326176
rect 93302 326136 93308 326148
rect 93360 326136 93366 326188
rect 93486 326176 93492 326188
rect 93447 326148 93492 326176
rect 93486 326136 93492 326148
rect 93544 326176 93550 326188
rect 117774 326176 117780 326188
rect 93544 326148 117780 326176
rect 93544 326136 93550 326148
rect 117774 326136 117780 326148
rect 117832 326136 117838 326188
rect 91557 326043 91615 326049
rect 91557 326009 91569 326043
rect 91603 326040 91615 326043
rect 91603 326012 103514 326040
rect 91603 326009 91615 326012
rect 91557 326003 91615 326009
rect 93673 325975 93731 325981
rect 93673 325941 93685 325975
rect 93719 325972 93731 325975
rect 103486 325972 103514 326012
rect 483014 325972 483020 325984
rect 93719 325944 93900 325972
rect 103486 325944 483020 325972
rect 93719 325941 93731 325944
rect 93673 325935 93731 325941
rect 93872 325768 93900 325944
rect 483014 325932 483020 325944
rect 483072 325932 483078 325984
rect 360838 325768 360844 325780
rect 93872 325740 360844 325768
rect 360838 325728 360844 325740
rect 360896 325728 360902 325780
rect 4706 325524 4712 325576
rect 4764 325564 4770 325576
rect 450541 325567 450599 325573
rect 450541 325564 450553 325567
rect 4764 325536 450553 325564
rect 4764 325524 4770 325536
rect 450541 325533 450553 325536
rect 450587 325533 450599 325567
rect 450541 325527 450599 325533
rect 331582 325088 331588 325100
rect 331495 325060 331588 325088
rect 331582 325048 331588 325060
rect 331640 325048 331646 325100
rect 331766 325048 331772 325100
rect 331824 325088 331830 325100
rect 385218 325088 385224 325100
rect 331824 325060 385224 325088
rect 331824 325048 331830 325060
rect 385218 325048 385224 325060
rect 385276 325048 385282 325100
rect 282270 325020 282276 325032
rect 282231 324992 282276 325020
rect 282270 324980 282276 324992
rect 282328 324980 282334 325032
rect 331600 325020 331628 325048
rect 385034 325020 385040 325032
rect 331600 324992 385040 325020
rect 385034 324980 385040 324992
rect 385092 324980 385098 325032
rect 277366 324924 287054 324952
rect 9214 324844 9220 324896
rect 9272 324884 9278 324896
rect 277366 324884 277394 324924
rect 9272 324856 277394 324884
rect 287026 324884 287054 324924
rect 331861 324887 331919 324893
rect 331861 324884 331873 324887
rect 287026 324856 331873 324884
rect 9272 324844 9278 324856
rect 331861 324853 331873 324856
rect 331907 324884 331919 324887
rect 423858 324884 423864 324896
rect 331907 324856 423864 324884
rect 331907 324853 331919 324856
rect 331861 324847 331919 324853
rect 423858 324844 423864 324856
rect 423916 324844 423922 324896
rect 400030 322872 400036 322924
rect 400088 322912 400094 322924
rect 495434 322912 495440 322924
rect 400088 322884 495440 322912
rect 400088 322872 400094 322884
rect 495434 322872 495440 322884
rect 495492 322872 495498 322924
rect 348418 322708 348424 322720
rect 348379 322680 348424 322708
rect 348418 322668 348424 322680
rect 348476 322668 348482 322720
rect 3602 321580 3608 321632
rect 3660 321620 3666 321632
rect 314470 321620 314476 321632
rect 3660 321592 314476 321620
rect 3660 321580 3666 321592
rect 314470 321580 314476 321592
rect 314528 321580 314534 321632
rect 401502 320152 401508 320204
rect 401560 320192 401566 320204
rect 465445 320195 465503 320201
rect 465445 320192 465457 320195
rect 401560 320164 465457 320192
rect 401560 320152 401566 320164
rect 465445 320161 465457 320164
rect 465491 320161 465503 320195
rect 465445 320155 465503 320161
rect 78953 319447 79011 319453
rect 78953 319413 78965 319447
rect 78999 319444 79011 319447
rect 313826 319444 313832 319456
rect 78999 319416 313832 319444
rect 78999 319413 79011 319416
rect 78953 319407 79011 319413
rect 313826 319404 313832 319416
rect 313884 319404 313890 319456
rect 342254 319104 342260 319116
rect 342215 319076 342260 319104
rect 342254 319064 342260 319076
rect 342312 319104 342318 319116
rect 342530 319104 342536 319116
rect 342312 319076 342536 319104
rect 342312 319064 342318 319076
rect 342530 319064 342536 319076
rect 342588 319064 342594 319116
rect 341990 318971 342048 318977
rect 341990 318937 342002 318971
rect 342036 318937 342048 318971
rect 341990 318931 342048 318937
rect 340877 318903 340935 318909
rect 340877 318869 340889 318903
rect 340923 318900 340935 318903
rect 340966 318900 340972 318912
rect 340923 318872 340972 318900
rect 340923 318869 340935 318872
rect 340877 318863 340935 318869
rect 340966 318860 340972 318872
rect 341024 318860 341030 318912
rect 341996 318900 342024 318931
rect 342070 318900 342076 318912
rect 341996 318872 342076 318900
rect 342070 318860 342076 318872
rect 342128 318860 342134 318912
rect 182082 317404 182088 317416
rect 182043 317376 182088 317404
rect 182082 317364 182088 317376
rect 182140 317364 182146 317416
rect 11698 317228 11704 317280
rect 11756 317268 11762 317280
rect 21269 317271 21327 317277
rect 21269 317268 21281 317271
rect 11756 317240 21281 317268
rect 11756 317228 11762 317240
rect 21269 317237 21281 317240
rect 21315 317237 21327 317271
rect 21269 317231 21327 317237
rect 481818 314344 481824 314356
rect 481779 314316 481824 314344
rect 481818 314304 481824 314316
rect 481876 314304 481882 314356
rect 481726 314208 481732 314220
rect 481687 314180 481732 314208
rect 481726 314168 481732 314180
rect 481784 314168 481790 314220
rect 64782 313216 64788 313268
rect 64840 313256 64846 313268
rect 495434 313256 495440 313268
rect 64840 313228 495440 313256
rect 64840 313216 64846 313228
rect 495434 313216 495440 313228
rect 495492 313216 495498 313268
rect 183373 312171 183431 312177
rect 183373 312168 183385 312171
rect 180766 312140 183385 312168
rect 7558 311856 7564 311908
rect 7616 311896 7622 311908
rect 180766 311896 180794 312140
rect 183373 312137 183385 312140
rect 183419 312168 183431 312171
rect 183419 312140 190454 312168
rect 183419 312137 183431 312140
rect 183373 312131 183431 312137
rect 184474 312060 184480 312112
rect 184532 312109 184538 312112
rect 184532 312100 184544 312109
rect 190426 312100 190454 312140
rect 412358 312100 412364 312112
rect 184532 312072 184577 312100
rect 190426 312072 412364 312100
rect 184532 312063 184544 312072
rect 184532 312060 184538 312063
rect 412358 312060 412364 312072
rect 412416 312060 412422 312112
rect 184753 311967 184811 311973
rect 184753 311933 184765 311967
rect 184799 311964 184811 311967
rect 243078 311964 243084 311976
rect 184799 311936 243084 311964
rect 184799 311933 184811 311936
rect 184753 311927 184811 311933
rect 243078 311924 243084 311936
rect 243136 311924 243142 311976
rect 7616 311868 180794 311896
rect 7616 311856 7622 311868
rect 23382 310700 23388 310752
rect 23440 310740 23446 310752
rect 403345 310743 403403 310749
rect 403345 310740 403357 310743
rect 23440 310712 403357 310740
rect 23440 310700 23446 310712
rect 403345 310709 403357 310712
rect 403391 310709 403403 310743
rect 403345 310703 403403 310709
rect 426710 308728 426716 308780
rect 426768 308768 426774 308780
rect 426805 308771 426863 308777
rect 426805 308768 426817 308771
rect 426768 308740 426817 308768
rect 426768 308728 426774 308740
rect 426805 308737 426817 308740
rect 426851 308737 426863 308771
rect 426805 308731 426863 308737
rect 426897 308771 426955 308777
rect 426897 308737 426909 308771
rect 426943 308768 426955 308771
rect 426986 308768 426992 308780
rect 426943 308740 426992 308768
rect 426943 308737 426955 308740
rect 426897 308731 426955 308737
rect 426986 308728 426992 308740
rect 427044 308728 427050 308780
rect 426437 308703 426495 308709
rect 426437 308700 426449 308703
rect 412606 308672 426449 308700
rect 380894 308592 380900 308644
rect 380952 308632 380958 308644
rect 412606 308632 412634 308672
rect 426437 308669 426449 308672
rect 426483 308669 426495 308703
rect 426437 308663 426495 308669
rect 426529 308703 426587 308709
rect 426529 308669 426541 308703
rect 426575 308700 426587 308703
rect 445754 308700 445760 308712
rect 426575 308672 445760 308700
rect 426575 308669 426587 308672
rect 426529 308663 426587 308669
rect 445754 308660 445760 308672
rect 445812 308660 445818 308712
rect 427081 308635 427139 308641
rect 427081 308632 427093 308635
rect 380952 308604 412634 308632
rect 424704 308604 427093 308632
rect 380952 308592 380958 308604
rect 264606 308524 264612 308576
rect 264664 308564 264670 308576
rect 424704 308564 424732 308604
rect 427081 308601 427093 308604
rect 427127 308601 427139 308635
rect 427081 308595 427139 308601
rect 264664 308536 424732 308564
rect 426437 308567 426495 308573
rect 264664 308524 264670 308536
rect 426437 308533 426449 308567
rect 426483 308564 426495 308567
rect 426621 308567 426679 308573
rect 426621 308564 426633 308567
rect 426483 308536 426633 308564
rect 426483 308533 426495 308536
rect 426437 308527 426495 308533
rect 426621 308533 426633 308536
rect 426667 308533 426679 308567
rect 426621 308527 426679 308533
rect 445754 308388 445760 308440
rect 445812 308428 445818 308440
rect 462314 308428 462320 308440
rect 445812 308400 462320 308428
rect 445812 308388 445818 308400
rect 462314 308388 462320 308400
rect 462372 308388 462378 308440
rect 483014 307776 483020 307828
rect 483072 307816 483078 307828
rect 495434 307816 495440 307828
rect 483072 307788 495440 307816
rect 483072 307776 483078 307788
rect 495434 307776 495440 307788
rect 495492 307776 495498 307828
rect 140685 307139 140743 307145
rect 140685 307105 140697 307139
rect 140731 307136 140743 307139
rect 140774 307136 140780 307148
rect 140731 307108 140780 307136
rect 140731 307105 140743 307108
rect 140685 307099 140743 307105
rect 140774 307096 140780 307108
rect 140832 307136 140838 307148
rect 180794 307136 180800 307148
rect 140832 307108 180800 307136
rect 140832 307096 140838 307108
rect 180794 307096 180800 307108
rect 180852 307096 180858 307148
rect 140774 307000 140780 307012
rect 140735 306972 140780 307000
rect 140774 306960 140780 306972
rect 140832 306960 140838 307012
rect 140866 306892 140872 306944
rect 140924 306932 140930 306944
rect 141234 306932 141240 306944
rect 140924 306904 140969 306932
rect 141195 306904 141240 306932
rect 140924 306892 140930 306904
rect 141234 306892 141240 306904
rect 141292 306892 141298 306944
rect 187421 306391 187479 306397
rect 187421 306357 187433 306391
rect 187467 306388 187479 306391
rect 351178 306388 351184 306400
rect 187467 306360 351184 306388
rect 187467 306357 187479 306360
rect 187421 306351 187479 306357
rect 351178 306348 351184 306360
rect 351236 306348 351242 306400
rect 22094 306184 22100 306196
rect 22055 306156 22100 306184
rect 22094 306144 22100 306156
rect 22152 306144 22158 306196
rect 21468 306088 26234 306116
rect 21468 306057 21496 306088
rect 21453 306051 21511 306057
rect 21453 306017 21465 306051
rect 21499 306017 21511 306051
rect 21634 306048 21640 306060
rect 21595 306020 21640 306048
rect 21453 306011 21511 306017
rect 21634 306008 21640 306020
rect 21692 306008 21698 306060
rect 26206 306048 26234 306088
rect 71866 306048 71872 306060
rect 26206 306020 71872 306048
rect 71866 306008 71872 306020
rect 71924 306008 71930 306060
rect 21542 305804 21548 305856
rect 21600 305844 21606 305856
rect 21729 305847 21787 305853
rect 21729 305844 21741 305847
rect 21600 305816 21741 305844
rect 21600 305804 21606 305816
rect 21729 305813 21741 305816
rect 21775 305813 21787 305847
rect 21729 305807 21787 305813
rect 49881 304895 49939 304901
rect 49881 304861 49893 304895
rect 49927 304892 49939 304895
rect 50065 304895 50123 304901
rect 50065 304892 50077 304895
rect 49927 304864 50077 304892
rect 49927 304861 49939 304864
rect 49881 304855 49939 304861
rect 50065 304861 50077 304864
rect 50111 304892 50123 304895
rect 61102 304892 61108 304904
rect 50111 304864 61108 304892
rect 50111 304861 50123 304864
rect 50065 304855 50123 304861
rect 61102 304852 61108 304864
rect 61160 304852 61166 304904
rect 11422 304784 11428 304836
rect 11480 304824 11486 304836
rect 50310 304827 50368 304833
rect 50310 304824 50322 304827
rect 11480 304796 50322 304824
rect 11480 304784 11486 304796
rect 50310 304793 50322 304796
rect 50356 304793 50368 304827
rect 50310 304787 50368 304793
rect 3878 304716 3884 304768
rect 3936 304756 3942 304768
rect 5810 304756 5816 304768
rect 3936 304728 5816 304756
rect 3936 304716 3942 304728
rect 5810 304716 5816 304728
rect 5868 304716 5874 304768
rect 51442 304756 51448 304768
rect 51355 304728 51448 304756
rect 51442 304716 51448 304728
rect 51500 304756 51506 304768
rect 153378 304756 153384 304768
rect 51500 304728 153384 304756
rect 51500 304716 51506 304728
rect 153378 304716 153384 304728
rect 153436 304716 153442 304768
rect 5902 304552 5908 304564
rect 5828 304524 5908 304552
rect 5828 304493 5856 304524
rect 5902 304512 5908 304524
rect 5960 304512 5966 304564
rect 5822 304487 5880 304493
rect 5822 304453 5834 304487
rect 5868 304453 5880 304487
rect 5822 304447 5880 304453
rect 6089 304351 6147 304357
rect 6089 304317 6101 304351
rect 6135 304348 6147 304351
rect 49881 304351 49939 304357
rect 49881 304348 49893 304351
rect 6135 304320 49893 304348
rect 6135 304317 6147 304320
rect 6089 304311 6147 304317
rect 49881 304317 49893 304320
rect 49927 304317 49939 304351
rect 49881 304311 49939 304317
rect 4706 304212 4712 304224
rect 4667 304184 4712 304212
rect 4706 304172 4712 304184
rect 4764 304212 4770 304224
rect 495618 304212 495624 304224
rect 4764 304184 495624 304212
rect 4764 304172 4770 304184
rect 495618 304172 495624 304184
rect 495676 304172 495682 304224
rect 4154 303084 4160 303136
rect 4212 303124 4218 303136
rect 325789 303127 325847 303133
rect 325789 303124 325801 303127
rect 4212 303096 325801 303124
rect 4212 303084 4218 303096
rect 325789 303093 325801 303096
rect 325835 303093 325847 303127
rect 325789 303087 325847 303093
rect 262493 301631 262551 301637
rect 262493 301597 262505 301631
rect 262539 301628 262551 301631
rect 263594 301628 263600 301640
rect 262539 301600 263600 301628
rect 262539 301597 262551 301600
rect 262493 301591 262551 301597
rect 263594 301588 263600 301600
rect 263652 301588 263658 301640
rect 262226 301563 262284 301569
rect 262226 301529 262238 301563
rect 262272 301529 262284 301563
rect 262226 301523 262284 301529
rect 261110 301492 261116 301504
rect 261071 301464 261116 301492
rect 261110 301452 261116 301464
rect 261168 301452 261174 301504
rect 262232 301492 262260 301523
rect 262306 301492 262312 301504
rect 262232 301464 262312 301492
rect 262306 301452 262312 301464
rect 262364 301452 262370 301504
rect 344738 301452 344744 301504
rect 344796 301492 344802 301504
rect 483750 301492 483756 301504
rect 344796 301464 483756 301492
rect 344796 301452 344802 301464
rect 483750 301452 483756 301464
rect 483808 301452 483814 301504
rect 341061 301155 341119 301161
rect 341061 301121 341073 301155
rect 341107 301152 341119 301155
rect 344738 301152 344744 301164
rect 341107 301124 344744 301152
rect 341107 301121 341119 301124
rect 341061 301115 341119 301121
rect 344738 301112 344744 301124
rect 344796 301112 344802 301164
rect 201954 301044 201960 301096
rect 202012 301084 202018 301096
rect 340877 301087 340935 301093
rect 340877 301084 340889 301087
rect 202012 301056 340889 301084
rect 202012 301044 202018 301056
rect 340877 301053 340889 301056
rect 340923 301053 340935 301087
rect 340877 301047 340935 301053
rect 193858 300908 193864 300960
rect 193916 300948 193922 300960
rect 341245 300951 341303 300957
rect 341245 300948 341257 300951
rect 193916 300920 341257 300948
rect 193916 300908 193922 300920
rect 341245 300917 341257 300920
rect 341291 300917 341303 300951
rect 341245 300911 341303 300917
rect 7834 300092 7840 300144
rect 7892 300132 7898 300144
rect 495434 300132 495440 300144
rect 7892 300104 495440 300132
rect 7892 300092 7898 300104
rect 495434 300092 495440 300104
rect 495492 300092 495498 300144
rect 3878 298324 3884 298376
rect 3936 298364 3942 298376
rect 46477 298367 46535 298373
rect 46477 298364 46489 298367
rect 3936 298336 46489 298364
rect 3936 298324 3942 298336
rect 46477 298333 46489 298336
rect 46523 298333 46535 298367
rect 46477 298327 46535 298333
rect 204990 296188 204996 296200
rect 200086 296160 204996 296188
rect 131114 295944 131120 295996
rect 131172 295984 131178 295996
rect 132402 295984 132408 295996
rect 131172 295956 132408 295984
rect 131172 295944 131178 295956
rect 132402 295944 132408 295956
rect 132460 295984 132466 295996
rect 200086 295984 200114 296160
rect 204990 296148 204996 296160
rect 205048 296188 205054 296200
rect 414201 296191 414259 296197
rect 414201 296188 414213 296191
rect 205048 296160 414213 296188
rect 205048 296148 205054 296160
rect 414201 296157 414213 296160
rect 414247 296157 414259 296191
rect 414382 296188 414388 296200
rect 414343 296160 414388 296188
rect 414201 296151 414259 296157
rect 414382 296148 414388 296160
rect 414440 296148 414446 296200
rect 262306 296012 262312 296064
rect 262364 296052 262370 296064
rect 414569 296055 414627 296061
rect 414569 296052 414581 296055
rect 262364 296024 414581 296052
rect 262364 296012 262370 296024
rect 414569 296021 414581 296024
rect 414615 296021 414627 296055
rect 414569 296015 414627 296021
rect 132460 295956 200114 295984
rect 132460 295944 132466 295956
rect 112809 295851 112867 295857
rect 112809 295817 112821 295851
rect 112855 295848 112867 295851
rect 259086 295848 259092 295860
rect 112855 295820 259092 295848
rect 112855 295817 112867 295820
rect 112809 295811 112867 295817
rect 259086 295808 259092 295820
rect 259144 295808 259150 295860
rect 131114 295780 131120 295792
rect 111996 295752 131120 295780
rect 111996 295721 112024 295752
rect 131114 295740 131120 295752
rect 131172 295740 131178 295792
rect 111981 295715 112039 295721
rect 111981 295681 111993 295715
rect 112027 295681 112039 295715
rect 111981 295675 112039 295681
rect 8294 295604 8300 295656
rect 8352 295644 8358 295656
rect 111996 295644 112024 295675
rect 112162 295672 112168 295724
rect 112220 295712 112226 295724
rect 112530 295712 112536 295724
rect 112220 295684 112264 295712
rect 112491 295684 112536 295712
rect 112220 295672 112226 295684
rect 112530 295672 112536 295684
rect 112588 295712 112594 295724
rect 112588 295684 113174 295712
rect 112588 295672 112594 295684
rect 8352 295616 112024 295644
rect 112257 295647 112315 295653
rect 8352 295604 8358 295616
rect 112257 295613 112269 295647
rect 112303 295613 112315 295647
rect 112257 295607 112315 295613
rect 112349 295647 112407 295653
rect 112349 295613 112361 295647
rect 112395 295644 112407 295647
rect 112809 295647 112867 295653
rect 112809 295644 112821 295647
rect 112395 295616 112821 295644
rect 112395 295613 112407 295616
rect 112349 295607 112407 295613
rect 112809 295613 112821 295616
rect 112855 295613 112867 295647
rect 113146 295644 113174 295684
rect 114462 295672 114468 295724
rect 114520 295712 114526 295724
rect 496262 295712 496268 295724
rect 114520 295684 496268 295712
rect 114520 295672 114526 295684
rect 496262 295672 496268 295684
rect 496320 295672 496326 295724
rect 311066 295644 311072 295656
rect 113146 295616 311072 295644
rect 112809 295607 112867 295613
rect 112272 295576 112300 295607
rect 311066 295604 311072 295616
rect 311124 295604 311130 295656
rect 259454 295576 259460 295588
rect 112272 295548 259460 295576
rect 259454 295536 259460 295548
rect 259512 295536 259518 295588
rect 112625 295511 112683 295517
rect 112625 295477 112637 295511
rect 112671 295508 112683 295511
rect 392118 295508 392124 295520
rect 112671 295480 392124 295508
rect 112671 295477 112683 295480
rect 112625 295471 112683 295477
rect 392118 295468 392124 295480
rect 392176 295468 392182 295520
rect 244366 295264 244372 295316
rect 244424 295304 244430 295316
rect 495434 295304 495440 295316
rect 244424 295276 495440 295304
rect 244424 295264 244430 295276
rect 495434 295264 495440 295276
rect 495492 295264 495498 295316
rect 104529 294015 104587 294021
rect 104529 293981 104541 294015
rect 104575 294012 104587 294015
rect 324958 294012 324964 294024
rect 104575 293984 324964 294012
rect 104575 293981 104587 293984
rect 104529 293975 104587 293981
rect 324958 293972 324964 293984
rect 325016 293972 325022 294024
rect 274726 293332 274732 293344
rect 274687 293304 274732 293332
rect 274726 293292 274732 293304
rect 274784 293292 274790 293344
rect 84197 292927 84255 292933
rect 84197 292893 84209 292927
rect 84243 292924 84255 292927
rect 367094 292924 367100 292936
rect 84243 292896 367100 292924
rect 84243 292893 84255 292896
rect 84197 292887 84255 292893
rect 367094 292884 367100 292896
rect 367152 292884 367158 292936
rect 70578 292408 70584 292460
rect 70636 292448 70642 292460
rect 138181 292451 138239 292457
rect 138181 292448 138193 292451
rect 70636 292420 138193 292448
rect 70636 292408 70642 292420
rect 138181 292417 138193 292420
rect 138227 292417 138239 292451
rect 138181 292411 138239 292417
rect 137922 292380 137928 292392
rect 137883 292352 137928 292380
rect 137922 292340 137928 292352
rect 137980 292340 137986 292392
rect 139305 292247 139363 292253
rect 139305 292213 139317 292247
rect 139351 292244 139363 292247
rect 240134 292244 240140 292256
rect 139351 292216 240140 292244
rect 139351 292213 139363 292216
rect 139305 292207 139363 292213
rect 240134 292204 240140 292216
rect 240192 292204 240198 292256
rect 341168 291468 345014 291496
rect 340874 291360 340880 291372
rect 340835 291332 340880 291360
rect 340874 291320 340880 291332
rect 340932 291320 340938 291372
rect 341168 291360 341196 291468
rect 341246 291363 341304 291369
rect 341246 291360 341258 291363
rect 341168 291332 341258 291360
rect 341246 291329 341258 291332
rect 341292 291329 341304 291363
rect 341426 291360 341432 291372
rect 341387 291332 341432 291360
rect 341246 291323 341304 291329
rect 341426 291320 341432 291332
rect 341484 291320 341490 291372
rect 344986 291360 345014 291468
rect 393314 291360 393320 291372
rect 344986 291332 393320 291360
rect 393314 291320 393320 291332
rect 393372 291320 393378 291372
rect 341061 291295 341119 291301
rect 341061 291261 341073 291295
rect 341107 291261 341119 291295
rect 341061 291255 341119 291261
rect 341153 291295 341211 291301
rect 341153 291261 341165 291295
rect 341199 291292 341211 291295
rect 341334 291292 341340 291304
rect 341199 291264 341340 291292
rect 341199 291261 341211 291264
rect 341153 291255 341211 291261
rect 195054 291184 195060 291236
rect 195112 291224 195118 291236
rect 340693 291227 340751 291233
rect 340693 291224 340705 291227
rect 195112 291196 340705 291224
rect 195112 291184 195118 291196
rect 340693 291193 340705 291196
rect 340739 291193 340751 291227
rect 341076 291224 341104 291255
rect 341334 291252 341340 291264
rect 341392 291252 341398 291304
rect 341242 291224 341248 291236
rect 341076 291196 341248 291224
rect 340693 291187 340751 291193
rect 341242 291184 341248 291196
rect 341300 291184 341306 291236
rect 3602 289824 3608 289876
rect 3660 289864 3666 289876
rect 312446 289864 312452 289876
rect 3660 289836 312452 289864
rect 3660 289824 3666 289836
rect 312446 289824 312452 289836
rect 312504 289824 312510 289876
rect 92934 288096 92940 288108
rect 92895 288068 92940 288096
rect 92934 288056 92940 288068
rect 92992 288056 92998 288108
rect 93118 288096 93124 288108
rect 93079 288068 93124 288096
rect 93118 288056 93124 288068
rect 93176 288056 93182 288108
rect 255682 288096 255688 288108
rect 93826 288068 255688 288096
rect 92952 288028 92980 288056
rect 93826 288028 93854 288068
rect 255682 288056 255688 288068
rect 255740 288056 255746 288108
rect 92952 288000 93854 288028
rect 59630 287852 59636 287904
rect 59688 287892 59694 287904
rect 92753 287895 92811 287901
rect 92753 287892 92765 287895
rect 59688 287864 92765 287892
rect 59688 287852 59694 287864
rect 92753 287861 92765 287864
rect 92799 287861 92811 287895
rect 92753 287855 92811 287861
rect 273622 287008 273628 287020
rect 273583 286980 273628 287008
rect 273622 286968 273628 286980
rect 273680 286968 273686 287020
rect 273806 287008 273812 287020
rect 273767 286980 273812 287008
rect 273806 286968 273812 286980
rect 273864 286968 273870 287020
rect 108298 286900 108304 286952
rect 108356 286940 108362 286952
rect 495434 286940 495440 286952
rect 108356 286912 495440 286940
rect 108356 286900 108362 286912
rect 495434 286900 495440 286912
rect 495492 286900 495498 286952
rect 273990 286872 273996 286884
rect 273951 286844 273996 286872
rect 273990 286832 273996 286844
rect 274048 286832 274054 286884
rect 244458 283880 244464 283892
rect 244419 283852 244464 283880
rect 244458 283840 244464 283852
rect 244516 283840 244522 283892
rect 134334 283704 134340 283756
rect 134392 283744 134398 283756
rect 243337 283747 243395 283753
rect 243337 283744 243349 283747
rect 134392 283716 243349 283744
rect 134392 283704 134398 283716
rect 243337 283713 243349 283716
rect 243383 283713 243395 283747
rect 263594 283744 263600 283756
rect 243337 283707 243395 283713
rect 248386 283716 263600 283744
rect 243078 283676 243084 283688
rect 242991 283648 243084 283676
rect 243078 283636 243084 283648
rect 243136 283636 243142 283688
rect 243096 283540 243124 283636
rect 248386 283608 248414 283716
rect 263594 283704 263600 283716
rect 263652 283704 263658 283756
rect 297545 283747 297603 283753
rect 297545 283713 297557 283747
rect 297591 283744 297603 283747
rect 297634 283744 297640 283756
rect 297591 283716 297640 283744
rect 297591 283713 297603 283716
rect 297545 283707 297603 283713
rect 297634 283704 297640 283716
rect 297692 283704 297698 283756
rect 296898 283636 296904 283688
rect 296956 283676 296962 283688
rect 297269 283679 297327 283685
rect 297269 283676 297281 283679
rect 296956 283648 297281 283676
rect 296956 283636 296962 283648
rect 297269 283645 297281 283648
rect 297315 283645 297327 283679
rect 297269 283639 297327 283645
rect 244016 283580 248414 283608
rect 244016 283540 244044 283580
rect 243096 283512 244044 283540
rect 244458 283500 244464 283552
rect 244516 283540 244522 283552
rect 257154 283540 257160 283552
rect 244516 283512 257160 283540
rect 244516 283500 244522 283512
rect 257154 283500 257160 283512
rect 257212 283500 257218 283552
rect 296070 283336 296076 283348
rect 296031 283308 296076 283336
rect 296070 283296 296076 283308
rect 296128 283296 296134 283348
rect 483014 283336 483020 283348
rect 482975 283308 483020 283336
rect 483014 283296 483020 283308
rect 483072 283296 483078 283348
rect 297634 283200 297640 283212
rect 297595 283172 297640 283200
rect 297634 283160 297640 283172
rect 297692 283160 297698 283212
rect 296257 283135 296315 283141
rect 296257 283101 296269 283135
rect 296303 283101 296315 283135
rect 296257 283095 296315 283101
rect 296272 283064 296300 283095
rect 296714 283092 296720 283144
rect 296772 283132 296778 283144
rect 296772 283104 296817 283132
rect 296772 283092 296778 283104
rect 296898 283064 296904 283076
rect 296272 283036 296904 283064
rect 296898 283024 296904 283036
rect 296956 283024 296962 283076
rect 296257 282795 296315 282801
rect 296257 282761 296269 282795
rect 296303 282792 296315 282795
rect 296714 282792 296720 282804
rect 296303 282764 296720 282792
rect 296303 282761 296315 282764
rect 296257 282755 296315 282761
rect 296714 282752 296720 282764
rect 296772 282752 296778 282804
rect 296070 282656 296076 282668
rect 296031 282628 296076 282656
rect 296070 282616 296076 282628
rect 296128 282616 296134 282668
rect 296898 282656 296904 282668
rect 296859 282628 296904 282656
rect 296898 282616 296904 282628
rect 296956 282616 296962 282668
rect 297913 282591 297971 282597
rect 297913 282557 297925 282591
rect 297959 282588 297971 282591
rect 321462 282588 321468 282600
rect 297959 282560 321468 282588
rect 297959 282557 297971 282560
rect 297913 282551 297971 282557
rect 321462 282548 321468 282560
rect 321520 282548 321526 282600
rect 296070 282480 296076 282532
rect 296128 282520 296134 282532
rect 296128 282492 335354 282520
rect 296128 282480 296134 282492
rect 335326 282180 335354 282492
rect 337746 282180 337752 282192
rect 335326 282152 337752 282180
rect 337746 282140 337752 282152
rect 337804 282180 337810 282192
rect 367554 282180 367560 282192
rect 337804 282152 367560 282180
rect 337804 282140 337810 282152
rect 367554 282140 367560 282152
rect 367612 282140 367618 282192
rect 16853 282047 16911 282053
rect 16853 282013 16865 282047
rect 16899 282044 16911 282047
rect 369210 282044 369216 282056
rect 16899 282016 369216 282044
rect 16899 282013 16911 282016
rect 16853 282007 16911 282013
rect 369210 282004 369216 282016
rect 369268 282004 369274 282056
rect 227898 281528 227904 281580
rect 227956 281568 227962 281580
rect 495434 281568 495440 281580
rect 227956 281540 495440 281568
rect 227956 281528 227962 281540
rect 495434 281528 495440 281540
rect 495492 281528 495498 281580
rect 5626 281324 5632 281376
rect 5684 281364 5690 281376
rect 84565 281367 84623 281373
rect 84565 281364 84577 281367
rect 5684 281336 84577 281364
rect 5684 281324 5690 281336
rect 84565 281333 84577 281336
rect 84611 281333 84623 281367
rect 84565 281327 84623 281333
rect 329742 280480 329748 280492
rect 329655 280452 329748 280480
rect 329742 280440 329748 280452
rect 329800 280480 329806 280492
rect 406286 280480 406292 280492
rect 329800 280452 406292 280480
rect 329800 280440 329806 280452
rect 406286 280440 406292 280452
rect 406344 280440 406350 280492
rect 135898 280236 135904 280288
rect 135956 280276 135962 280288
rect 329653 280279 329711 280285
rect 329653 280276 329665 280279
rect 135956 280248 329665 280276
rect 135956 280236 135962 280248
rect 329653 280245 329665 280248
rect 329699 280245 329711 280279
rect 329653 280239 329711 280245
rect 264606 279469 264612 279472
rect 264600 279460 264612 279469
rect 264567 279432 264612 279460
rect 264600 279423 264612 279432
rect 264606 279420 264612 279423
rect 264664 279420 264670 279472
rect 263594 279352 263600 279404
rect 263652 279392 263658 279404
rect 264333 279395 264391 279401
rect 264333 279392 264345 279395
rect 263652 279364 264345 279392
rect 263652 279352 263658 279364
rect 264333 279361 264345 279364
rect 264379 279392 264391 279395
rect 266354 279392 266360 279404
rect 264379 279364 266360 279392
rect 264379 279361 264391 279364
rect 264333 279355 264391 279361
rect 266354 279352 266360 279364
rect 266412 279352 266418 279404
rect 265713 279191 265771 279197
rect 265713 279157 265725 279191
rect 265759 279188 265771 279191
rect 426894 279188 426900 279200
rect 265759 279160 426900 279188
rect 265759 279157 265771 279160
rect 265713 279151 265771 279157
rect 426894 279148 426900 279160
rect 426952 279148 426958 279200
rect 176930 277896 176936 277908
rect 176891 277868 176936 277896
rect 176930 277856 176936 277868
rect 176988 277856 176994 277908
rect 248690 276128 248696 276140
rect 248651 276100 248696 276128
rect 248690 276088 248696 276100
rect 248748 276088 248754 276140
rect 248598 276060 248604 276072
rect 248559 276032 248604 276060
rect 248598 276020 248604 276032
rect 248656 276020 248662 276072
rect 158916 273992 161474 274020
rect 158916 273964 158944 273992
rect 125870 273912 125876 273964
rect 125928 273952 125934 273964
rect 158717 273955 158775 273961
rect 158717 273952 158729 273955
rect 125928 273924 158729 273952
rect 125928 273912 125934 273924
rect 158717 273921 158729 273924
rect 158763 273921 158775 273955
rect 158898 273952 158904 273964
rect 158859 273924 158904 273952
rect 158717 273915 158775 273921
rect 158898 273912 158904 273924
rect 158956 273912 158962 273964
rect 159082 273952 159088 273964
rect 159043 273924 159088 273952
rect 159082 273912 159088 273924
rect 159140 273912 159146 273964
rect 159266 273952 159272 273964
rect 159227 273924 159272 273952
rect 159266 273912 159272 273924
rect 159324 273912 159330 273964
rect 161446 273952 161474 273992
rect 248230 273952 248236 273964
rect 161446 273924 248236 273952
rect 248230 273912 248236 273924
rect 248288 273952 248294 273964
rect 402790 273952 402796 273964
rect 248288 273924 402796 273952
rect 248288 273912 248294 273924
rect 402790 273912 402796 273924
rect 402848 273912 402854 273964
rect 158990 273884 158996 273896
rect 158951 273856 158996 273884
rect 158990 273844 158996 273856
rect 159048 273844 159054 273896
rect 159100 273884 159128 273912
rect 248598 273884 248604 273896
rect 159100 273856 248604 273884
rect 248598 273844 248604 273856
rect 248656 273844 248662 273896
rect 89162 273708 89168 273760
rect 89220 273748 89226 273760
rect 159361 273751 159419 273757
rect 159361 273748 159373 273751
rect 89220 273720 159373 273748
rect 89220 273708 89226 273720
rect 159361 273717 159373 273720
rect 159407 273717 159419 273751
rect 159361 273711 159419 273717
rect 3234 273300 3240 273352
rect 3292 273340 3298 273352
rect 229097 273343 229155 273349
rect 229097 273340 229109 273343
rect 3292 273312 229109 273340
rect 3292 273300 3298 273312
rect 229097 273309 229109 273312
rect 229143 273309 229155 273343
rect 229097 273303 229155 273309
rect 3602 273164 3608 273216
rect 3660 273204 3666 273216
rect 207106 273204 207112 273216
rect 3660 273176 207112 273204
rect 3660 273164 3666 273176
rect 207106 273164 207112 273176
rect 207164 273164 207170 273216
rect 420546 272660 420552 272672
rect 420507 272632 420552 272660
rect 420546 272620 420552 272632
rect 420604 272620 420610 272672
rect 373074 271328 373080 271380
rect 373132 271368 373138 271380
rect 375466 271368 375472 271380
rect 373132 271340 375472 271368
rect 373132 271328 373138 271340
rect 375466 271328 375472 271340
rect 375524 271328 375530 271380
rect 373261 271303 373319 271309
rect 373261 271269 373273 271303
rect 373307 271300 373319 271303
rect 373307 271272 373764 271300
rect 373307 271269 373319 271272
rect 373261 271263 373319 271269
rect 221458 271124 221464 271176
rect 221516 271164 221522 271176
rect 310698 271164 310704 271176
rect 221516 271136 310704 271164
rect 221516 271124 221522 271136
rect 310698 271124 310704 271136
rect 310756 271124 310762 271176
rect 373074 271164 373080 271176
rect 373035 271136 373080 271164
rect 373074 271124 373080 271136
rect 373132 271124 373138 271176
rect 373736 271173 373764 271272
rect 373721 271167 373779 271173
rect 373721 271133 373733 271167
rect 373767 271133 373779 271167
rect 373721 271127 373779 271133
rect 374917 271099 374975 271105
rect 374917 271065 374929 271099
rect 374963 271096 374975 271099
rect 375285 271099 375343 271105
rect 375285 271096 375297 271099
rect 374963 271068 375297 271096
rect 374963 271065 374975 271068
rect 374917 271059 374975 271065
rect 375285 271065 375297 271068
rect 375331 271096 375343 271099
rect 406378 271096 406384 271108
rect 375331 271068 406384 271096
rect 375331 271065 375343 271068
rect 375285 271059 375343 271065
rect 406378 271056 406384 271068
rect 406436 271056 406442 271108
rect 373810 270824 373816 270836
rect 373771 270796 373816 270824
rect 373810 270784 373816 270796
rect 373868 270784 373874 270836
rect 374273 270691 374331 270697
rect 374273 270657 374285 270691
rect 374319 270688 374331 270691
rect 375285 270691 375343 270697
rect 375285 270688 375297 270691
rect 374319 270660 375297 270688
rect 374319 270657 374331 270660
rect 374273 270651 374331 270657
rect 375285 270657 375297 270660
rect 375331 270657 375343 270691
rect 375285 270651 375343 270657
rect 92290 270280 92296 270292
rect 92251 270252 92296 270280
rect 92290 270240 92296 270252
rect 92348 270240 92354 270292
rect 92477 270079 92535 270085
rect 92477 270045 92489 270079
rect 92523 270076 92535 270079
rect 296070 270076 296076 270088
rect 92523 270048 296076 270076
rect 92523 270045 92535 270048
rect 92477 270039 92535 270045
rect 296070 270036 296076 270048
rect 296128 270036 296134 270088
rect 92290 269900 92296 269952
rect 92348 269940 92354 269952
rect 298830 269940 298836 269952
rect 92348 269912 298836 269940
rect 92348 269900 92354 269912
rect 298830 269900 298836 269912
rect 298888 269900 298894 269952
rect 141234 267860 141240 267912
rect 141292 267900 141298 267912
rect 228729 267903 228787 267909
rect 228729 267900 228741 267903
rect 141292 267872 228741 267900
rect 141292 267860 141298 267872
rect 228729 267869 228741 267872
rect 228775 267869 228787 267903
rect 228729 267863 228787 267869
rect 228910 267860 228916 267912
rect 228968 267900 228974 267912
rect 310238 267900 310244 267912
rect 228968 267872 310244 267900
rect 228968 267860 228974 267872
rect 310238 267860 310244 267872
rect 310296 267860 310302 267912
rect 219406 267804 238754 267832
rect 3602 267724 3608 267776
rect 3660 267764 3666 267776
rect 219406 267764 219434 267804
rect 3660 267736 219434 267764
rect 3660 267724 3666 267736
rect 229094 267724 229100 267776
rect 229152 267764 229158 267776
rect 238726 267764 238754 267804
rect 252554 267764 252560 267776
rect 229152 267736 229197 267764
rect 238726 267736 252560 267764
rect 229152 267724 229158 267736
rect 252554 267724 252560 267736
rect 252612 267724 252618 267776
rect 315482 267724 315488 267776
rect 315540 267764 315546 267776
rect 495434 267764 495440 267776
rect 315540 267736 495440 267764
rect 315540 267724 315546 267736
rect 495434 267724 495440 267736
rect 495492 267724 495498 267776
rect 367278 266812 367284 266824
rect 367239 266784 367284 266812
rect 367278 266772 367284 266784
rect 367336 266772 367342 266824
rect 367462 266812 367468 266824
rect 367423 266784 367468 266812
rect 367462 266772 367468 266784
rect 367520 266772 367526 266824
rect 486970 266812 486976 266824
rect 486931 266784 486976 266812
rect 486970 266772 486976 266784
rect 487028 266772 487034 266824
rect 299382 266704 299388 266756
rect 299440 266744 299446 266756
rect 486706 266747 486764 266753
rect 486706 266744 486718 266747
rect 299440 266716 486718 266744
rect 299440 266704 299446 266716
rect 486706 266713 486718 266716
rect 486752 266713 486764 266747
rect 486706 266707 486764 266713
rect 53926 266636 53932 266688
rect 53984 266676 53990 266688
rect 367097 266679 367155 266685
rect 367097 266676 367109 266679
rect 53984 266648 367109 266676
rect 53984 266636 53990 266648
rect 367097 266645 367109 266648
rect 367143 266645 367155 266679
rect 485590 266676 485596 266688
rect 485551 266648 485596 266676
rect 367097 266639 367155 266645
rect 485590 266636 485596 266648
rect 485648 266636 485654 266688
rect 36354 266336 36360 266348
rect 36315 266308 36360 266336
rect 36354 266296 36360 266308
rect 36412 266296 36418 266348
rect 86862 265752 86868 265804
rect 86920 265792 86926 265804
rect 353389 265795 353447 265801
rect 353389 265792 353401 265795
rect 86920 265764 353401 265792
rect 86920 265752 86926 265764
rect 353389 265761 353401 265764
rect 353435 265761 353447 265795
rect 353389 265755 353447 265761
rect 6730 265684 6736 265736
rect 6788 265724 6794 265736
rect 442261 265727 442319 265733
rect 442261 265724 442273 265727
rect 6788 265696 335354 265724
rect 6788 265684 6794 265696
rect 335326 265656 335354 265696
rect 354646 265696 442273 265724
rect 354646 265656 354674 265696
rect 442261 265693 442273 265696
rect 442307 265693 442319 265727
rect 442261 265687 442319 265693
rect 335326 265628 354674 265656
rect 78122 264169 78128 264172
rect 78116 264123 78128 264169
rect 78180 264160 78186 264172
rect 78180 264132 78216 264160
rect 78122 264120 78128 264123
rect 78180 264120 78186 264132
rect 77846 264092 77852 264104
rect 77807 264064 77852 264092
rect 77846 264052 77852 264064
rect 77904 264052 77910 264104
rect 84166 263996 103514 264024
rect 9030 263916 9036 263968
rect 9088 263956 9094 263968
rect 79226 263956 79232 263968
rect 9088 263928 79232 263956
rect 9088 263916 9094 263928
rect 79226 263916 79232 263928
rect 79284 263956 79290 263968
rect 84166 263956 84194 263996
rect 98730 263956 98736 263968
rect 79284 263928 84194 263956
rect 98691 263928 98736 263956
rect 79284 263916 79290 263928
rect 98730 263916 98736 263928
rect 98788 263916 98794 263968
rect 103486 263956 103514 263996
rect 331398 263956 331404 263968
rect 103486 263928 331404 263956
rect 331398 263916 331404 263928
rect 331456 263916 331462 263968
rect 207198 262556 207204 262608
rect 207256 262596 207262 262608
rect 207385 262599 207443 262605
rect 207385 262596 207397 262599
rect 207256 262568 207397 262596
rect 207256 262556 207262 262568
rect 207385 262565 207397 262568
rect 207431 262565 207443 262599
rect 207385 262559 207443 262565
rect 207014 262420 207020 262472
rect 207072 262460 207078 262472
rect 207109 262463 207167 262469
rect 207109 262460 207121 262463
rect 207072 262432 207121 262460
rect 207072 262420 207078 262432
rect 207109 262429 207121 262432
rect 207155 262429 207167 262463
rect 207382 262460 207388 262472
rect 207343 262432 207388 262460
rect 207109 262423 207167 262429
rect 207382 262420 207388 262432
rect 207440 262460 207446 262472
rect 402974 262460 402980 262472
rect 207440 262432 402980 262460
rect 207440 262420 207446 262432
rect 402974 262420 402980 262432
rect 403032 262420 403038 262472
rect 130470 261264 130476 261316
rect 130528 261304 130534 261316
rect 158806 261304 158812 261316
rect 130528 261276 158812 261304
rect 130528 261264 130534 261276
rect 158806 261264 158812 261276
rect 158864 261264 158870 261316
rect 125778 261196 125784 261248
rect 125836 261236 125842 261248
rect 125836 261208 132494 261236
rect 125836 261196 125842 261208
rect 125870 261032 125876 261044
rect 125928 261041 125934 261044
rect 125839 261004 125876 261032
rect 125870 260992 125876 261004
rect 125928 260995 125939 261041
rect 126057 261035 126115 261041
rect 126057 261001 126069 261035
rect 126103 261032 126115 261035
rect 132466 261032 132494 261208
rect 273806 261032 273812 261044
rect 126103 261004 129964 261032
rect 132466 261004 273812 261032
rect 126103 261001 126115 261004
rect 126057 260995 126115 261001
rect 125928 260992 125934 260995
rect 125505 260967 125563 260973
rect 125505 260933 125517 260967
rect 125551 260964 125563 260967
rect 129936 260964 129964 261004
rect 273806 260992 273812 261004
rect 273864 260992 273870 261044
rect 319806 260964 319812 260976
rect 125551 260936 129872 260964
rect 129936 260936 319812 260964
rect 125551 260933 125563 260936
rect 125505 260927 125563 260933
rect 125318 260896 125324 260908
rect 125279 260868 125324 260896
rect 125318 260856 125324 260868
rect 125376 260856 125382 260908
rect 125778 260905 125784 260908
rect 125597 260899 125655 260905
rect 125597 260865 125609 260899
rect 125643 260865 125655 260899
rect 125597 260859 125655 260865
rect 125741 260899 125784 260905
rect 125741 260865 125753 260899
rect 125741 260859 125784 260865
rect 125612 260828 125640 260859
rect 125778 260856 125784 260859
rect 125836 260856 125842 260908
rect 125870 260856 125876 260908
rect 125928 260896 125934 260908
rect 126057 260899 126115 260905
rect 126057 260896 126069 260899
rect 125928 260868 126069 260896
rect 125928 260856 125934 260868
rect 126057 260865 126069 260868
rect 126103 260865 126115 260899
rect 129844 260896 129872 260936
rect 319806 260924 319812 260936
rect 319864 260924 319870 260976
rect 131574 260896 131580 260908
rect 129844 260868 131580 260896
rect 126057 260859 126115 260865
rect 131574 260856 131580 260868
rect 131632 260896 131638 260908
rect 319898 260896 319904 260908
rect 131632 260868 319904 260896
rect 131632 260856 131638 260868
rect 319898 260856 319904 260868
rect 319956 260856 319962 260908
rect 125888 260828 125916 260856
rect 125612 260800 125916 260828
rect 317785 260287 317843 260293
rect 317785 260253 317797 260287
rect 317831 260284 317843 260287
rect 339954 260284 339960 260296
rect 317831 260256 339960 260284
rect 317831 260253 317843 260256
rect 317785 260247 317843 260253
rect 339954 260244 339960 260256
rect 340012 260244 340018 260296
rect 317690 260148 317696 260160
rect 317603 260120 317696 260148
rect 317690 260108 317696 260120
rect 317748 260148 317754 260160
rect 331214 260148 331220 260160
rect 317748 260120 331220 260148
rect 317748 260108 317754 260120
rect 331214 260108 331220 260120
rect 331272 260108 331278 260160
rect 180705 259267 180763 259273
rect 180705 259233 180717 259267
rect 180751 259264 180763 259267
rect 180794 259264 180800 259276
rect 180751 259236 180800 259264
rect 180751 259233 180763 259236
rect 180705 259227 180763 259233
rect 180794 259224 180800 259236
rect 180852 259264 180858 259276
rect 180978 259264 180984 259276
rect 180852 259236 180984 259264
rect 180852 259224 180858 259236
rect 180978 259224 180984 259236
rect 181036 259264 181042 259276
rect 232682 259264 232688 259276
rect 181036 259236 232688 259264
rect 181036 259224 181042 259236
rect 232682 259224 232688 259236
rect 232740 259224 232746 259276
rect 60001 259199 60059 259205
rect 60001 259165 60013 259199
rect 60047 259196 60059 259199
rect 268378 259196 268384 259208
rect 60047 259168 268384 259196
rect 60047 259165 60059 259168
rect 60001 259159 60059 259165
rect 268378 259156 268384 259168
rect 268436 259156 268442 259208
rect 180886 259128 180892 259140
rect 180847 259100 180892 259128
rect 180886 259088 180892 259100
rect 180944 259088 180950 259140
rect 180794 259020 180800 259072
rect 180852 259060 180858 259072
rect 181254 259060 181260 259072
rect 180852 259032 180897 259060
rect 181215 259032 181260 259060
rect 180852 259020 180858 259032
rect 181254 259020 181260 259032
rect 181312 259020 181318 259072
rect 347038 258068 347044 258120
rect 347096 258108 347102 258120
rect 495434 258108 495440 258120
rect 347096 258080 495440 258108
rect 347096 258068 347102 258080
rect 495434 258068 495440 258080
rect 495492 258068 495498 258120
rect 483750 257632 483756 257644
rect 483711 257604 483756 257632
rect 483750 257592 483756 257604
rect 483808 257592 483814 257644
rect 181254 257524 181260 257576
rect 181312 257564 181318 257576
rect 483569 257567 483627 257573
rect 483569 257564 483581 257567
rect 181312 257536 483581 257564
rect 181312 257524 181318 257536
rect 483569 257533 483581 257536
rect 483615 257533 483627 257567
rect 483569 257527 483627 257533
rect 321922 257388 321928 257440
rect 321980 257428 321986 257440
rect 483937 257431 483995 257437
rect 483937 257428 483949 257431
rect 321980 257400 483949 257428
rect 321980 257388 321986 257400
rect 483937 257397 483949 257400
rect 483983 257397 483995 257431
rect 483937 257391 483995 257397
rect 470502 257020 470508 257032
rect 470463 256992 470508 257020
rect 470502 256980 470508 256992
rect 470560 256980 470566 257032
rect 470594 256844 470600 256896
rect 470652 256884 470658 256896
rect 470652 256856 470697 256884
rect 470652 256844 470658 256856
rect 299382 256680 299388 256692
rect 299343 256652 299388 256680
rect 299382 256640 299388 256652
rect 299440 256640 299446 256692
rect 299109 256547 299167 256553
rect 299109 256544 299121 256547
rect 298664 256516 299121 256544
rect 298664 256408 298692 256516
rect 299109 256513 299121 256516
rect 299155 256513 299167 256547
rect 299109 256507 299167 256513
rect 299198 256504 299204 256556
rect 299256 256544 299262 256556
rect 485590 256544 485596 256556
rect 299256 256516 485596 256544
rect 299256 256504 299262 256516
rect 485590 256504 485596 256516
rect 485648 256504 485654 256556
rect 298830 256476 298836 256488
rect 298743 256448 298836 256476
rect 298830 256436 298836 256448
rect 298888 256476 298894 256488
rect 333974 256476 333980 256488
rect 298888 256448 333980 256476
rect 298888 256436 298894 256448
rect 333974 256436 333980 256448
rect 334032 256476 334038 256488
rect 334342 256476 334348 256488
rect 334032 256448 334348 256476
rect 334032 256436 334038 256448
rect 334342 256436 334348 256448
rect 334400 256436 334406 256488
rect 310422 256408 310428 256420
rect 298664 256380 310428 256408
rect 310422 256368 310428 256380
rect 310480 256368 310486 256420
rect 117590 256300 117596 256352
rect 117648 256340 117654 256352
rect 298925 256343 298983 256349
rect 298925 256340 298937 256343
rect 117648 256312 298937 256340
rect 117648 256300 117654 256312
rect 298925 256309 298937 256312
rect 298971 256309 298983 256343
rect 298925 256303 298983 256309
rect 333974 256028 333980 256080
rect 334032 256068 334038 256080
rect 371142 256068 371148 256080
rect 334032 256040 371148 256068
rect 334032 256028 334038 256040
rect 371142 256028 371148 256040
rect 371200 256028 371206 256080
rect 310054 255960 310060 256012
rect 310112 256000 310118 256012
rect 310422 256000 310428 256012
rect 310112 255972 310428 256000
rect 310112 255960 310118 255972
rect 310422 255960 310428 255972
rect 310480 256000 310486 256012
rect 334066 256000 334072 256012
rect 310480 255972 334072 256000
rect 310480 255960 310486 255972
rect 334066 255960 334072 255972
rect 334124 256000 334130 256012
rect 371418 256000 371424 256012
rect 334124 255972 371424 256000
rect 334124 255960 334130 255972
rect 371418 255960 371424 255972
rect 371476 255960 371482 256012
rect 263778 255212 263784 255264
rect 263836 255252 263842 255264
rect 381446 255252 381452 255264
rect 263836 255224 381452 255252
rect 263836 255212 263842 255224
rect 381446 255212 381452 255224
rect 381504 255212 381510 255264
rect 220538 254912 220544 254924
rect 220499 254884 220544 254912
rect 220538 254872 220544 254884
rect 220596 254872 220602 254924
rect 396626 254844 396632 254856
rect 396587 254816 396632 254844
rect 396626 254804 396632 254816
rect 396684 254804 396690 254856
rect 219802 254736 219808 254788
rect 219860 254776 219866 254788
rect 220274 254779 220332 254785
rect 220274 254776 220286 254779
rect 219860 254748 220286 254776
rect 219860 254736 219866 254748
rect 220274 254745 220286 254748
rect 220320 254745 220332 254779
rect 220274 254739 220332 254745
rect 219161 254711 219219 254717
rect 219161 254677 219173 254711
rect 219207 254708 219219 254711
rect 219250 254708 219256 254720
rect 219207 254680 219256 254708
rect 219207 254677 219219 254680
rect 219161 254671 219219 254677
rect 219250 254668 219256 254680
rect 219308 254708 219314 254720
rect 263778 254708 263784 254720
rect 219308 254680 263784 254708
rect 219308 254668 219314 254680
rect 263778 254668 263784 254680
rect 263836 254668 263842 254720
rect 349062 254124 349068 254176
rect 349120 254164 349126 254176
rect 380621 254167 380679 254173
rect 380621 254164 380633 254167
rect 349120 254136 380633 254164
rect 349120 254124 349126 254136
rect 380621 254133 380633 254136
rect 380667 254133 380679 254167
rect 380621 254127 380679 254133
rect 117590 252872 117596 252884
rect 117551 252844 117596 252872
rect 117590 252832 117596 252844
rect 117648 252832 117654 252884
rect 139029 252807 139087 252813
rect 139029 252804 139041 252807
rect 122806 252776 139041 252804
rect 3234 252696 3240 252748
rect 3292 252736 3298 252748
rect 122806 252736 122834 252776
rect 139029 252773 139041 252776
rect 139075 252773 139087 252807
rect 139029 252767 139087 252773
rect 3292 252708 122834 252736
rect 137296 252708 142154 252736
rect 3292 252696 3298 252708
rect 9306 252628 9312 252680
rect 9364 252668 9370 252680
rect 117774 252668 117780 252680
rect 9364 252640 117780 252668
rect 9364 252628 9370 252640
rect 117774 252628 117780 252640
rect 117832 252628 117838 252680
rect 117961 252671 118019 252677
rect 117961 252637 117973 252671
rect 118007 252668 118019 252671
rect 137296 252668 137324 252708
rect 118007 252640 137324 252668
rect 142126 252668 142154 252708
rect 414658 252668 414664 252680
rect 142126 252640 414664 252668
rect 118007 252637 118019 252640
rect 117961 252631 118019 252637
rect 414658 252628 414664 252640
rect 414716 252628 414722 252680
rect 117792 252600 117820 252628
rect 260650 252600 260656 252612
rect 117792 252572 260656 252600
rect 260650 252560 260656 252572
rect 260708 252560 260714 252612
rect 444006 252192 444012 252204
rect 443967 252164 444012 252192
rect 444006 252152 444012 252164
rect 444064 252152 444070 252204
rect 444098 252124 444104 252136
rect 444059 252096 444104 252124
rect 444098 252084 444104 252096
rect 444156 252084 444162 252136
rect 444190 252084 444196 252136
rect 444248 252124 444254 252136
rect 444248 252096 444293 252124
rect 444248 252084 444254 252096
rect 336090 251948 336096 252000
rect 336148 251988 336154 252000
rect 443641 251991 443699 251997
rect 443641 251988 443653 251991
rect 336148 251960 443653 251988
rect 336148 251948 336154 251960
rect 443641 251957 443653 251960
rect 443687 251957 443699 251991
rect 443641 251951 443699 251957
rect 274726 251132 274732 251184
rect 274784 251172 274790 251184
rect 495434 251172 495440 251184
rect 274784 251144 495440 251172
rect 274784 251132 274790 251144
rect 495434 251132 495440 251144
rect 495492 251132 495498 251184
rect 4614 251064 4620 251116
rect 4672 251104 4678 251116
rect 231193 251107 231251 251113
rect 231193 251104 231205 251107
rect 4672 251076 231205 251104
rect 4672 251064 4678 251076
rect 231193 251073 231205 251076
rect 231239 251073 231251 251107
rect 266354 251104 266360 251116
rect 231193 251067 231251 251073
rect 232240 251076 266360 251104
rect 230937 251039 230995 251045
rect 230937 251005 230949 251039
rect 230983 251005 230995 251039
rect 230937 250999 230995 251005
rect 230952 250900 230980 250999
rect 232240 250900 232268 251076
rect 266354 251064 266360 251076
rect 266412 251064 266418 251116
rect 232314 250928 232320 250980
rect 232372 250968 232378 250980
rect 232372 250940 238754 250968
rect 232372 250928 232378 250940
rect 230952 250872 232268 250900
rect 238726 250900 238754 250940
rect 254210 250900 254216 250912
rect 238726 250872 254216 250900
rect 254210 250860 254216 250872
rect 254268 250900 254274 250912
rect 257246 250900 257252 250912
rect 254268 250872 257252 250900
rect 254268 250860 254274 250872
rect 257246 250860 257252 250872
rect 257304 250860 257310 250912
rect 303154 250016 303160 250028
rect 303115 249988 303160 250016
rect 303154 249976 303160 249988
rect 303212 250016 303218 250028
rect 361574 250016 361580 250028
rect 303212 249988 361580 250016
rect 303212 249976 303218 249988
rect 361574 249976 361580 249988
rect 361632 249976 361638 250028
rect 12986 249772 12992 249824
rect 13044 249812 13050 249824
rect 302973 249815 303031 249821
rect 302973 249812 302985 249815
rect 13044 249784 302985 249812
rect 13044 249772 13050 249784
rect 302973 249781 302985 249784
rect 303019 249781 303031 249815
rect 302973 249775 303031 249781
rect 315114 248724 315120 248736
rect 315075 248696 315120 248724
rect 315114 248684 315120 248696
rect 315172 248684 315178 248736
rect 115201 244375 115259 244381
rect 115201 244341 115213 244375
rect 115247 244372 115259 244375
rect 311434 244372 311440 244384
rect 115247 244344 311440 244372
rect 115247 244341 115259 244344
rect 115201 244335 115259 244341
rect 311434 244332 311440 244344
rect 311492 244332 311498 244384
rect 315758 240904 315764 240916
rect 315719 240876 315764 240904
rect 315758 240864 315764 240876
rect 315816 240864 315822 240916
rect 468018 240904 468024 240916
rect 467979 240876 468024 240904
rect 468018 240864 468024 240876
rect 468076 240864 468082 240916
rect 467374 240632 467380 240644
rect 467335 240604 467380 240632
rect 467374 240592 467380 240604
rect 467432 240592 467438 240644
rect 467834 240632 467840 240644
rect 467795 240604 467840 240632
rect 467834 240592 467840 240604
rect 467892 240632 467898 240644
rect 496262 240632 496268 240644
rect 467892 240604 496268 240632
rect 467892 240592 467898 240604
rect 496262 240592 496268 240604
rect 496320 240592 496326 240644
rect 467650 240564 467656 240576
rect 467611 240536 467656 240564
rect 467650 240524 467656 240536
rect 467708 240524 467714 240576
rect 467742 240524 467748 240576
rect 467800 240564 467806 240576
rect 467800 240536 467845 240564
rect 467800 240524 467806 240536
rect 372614 238484 372620 238536
rect 372672 238524 372678 238536
rect 373074 238524 373080 238536
rect 372672 238496 373080 238524
rect 372672 238484 372678 238496
rect 373074 238484 373080 238496
rect 373132 238484 373138 238536
rect 20530 237572 20536 237584
rect 20491 237544 20536 237572
rect 20530 237532 20536 237544
rect 20588 237572 20594 237584
rect 430942 237572 430948 237584
rect 20588 237544 26234 237572
rect 430903 237544 430948 237572
rect 20588 237532 20594 237544
rect 26206 237504 26234 237544
rect 430942 237532 430948 237544
rect 431000 237532 431006 237584
rect 59446 237504 59452 237516
rect 26206 237476 59452 237504
rect 59446 237464 59452 237476
rect 59504 237464 59510 237516
rect 20349 237439 20407 237445
rect 20349 237405 20361 237439
rect 20395 237436 20407 237439
rect 372614 237436 372620 237448
rect 20395 237408 372620 237436
rect 20395 237405 20407 237408
rect 20349 237399 20407 237405
rect 372614 237396 372620 237408
rect 372672 237396 372678 237448
rect 430758 237436 430764 237448
rect 430719 237408 430764 237436
rect 430758 237396 430764 237408
rect 430816 237396 430822 237448
rect 430942 237396 430948 237448
rect 431000 237436 431006 237448
rect 435266 237436 435272 237448
rect 431000 237408 435272 237436
rect 431000 237396 431006 237408
rect 435266 237396 435272 237408
rect 435324 237396 435330 237448
rect 77846 236648 77852 236700
rect 77904 236688 77910 236700
rect 133230 236688 133236 236700
rect 77904 236660 133236 236688
rect 77904 236648 77910 236660
rect 133230 236648 133236 236660
rect 133288 236648 133294 236700
rect 5166 236308 5172 236360
rect 5224 236348 5230 236360
rect 61102 236348 61108 236360
rect 5224 236320 61108 236348
rect 5224 236308 5230 236320
rect 61102 236308 61108 236320
rect 61160 236348 61166 236360
rect 77846 236348 77852 236360
rect 61160 236320 77852 236348
rect 61160 236308 61166 236320
rect 77846 236308 77852 236320
rect 77904 236308 77910 236360
rect 342530 236348 342536 236360
rect 342491 236320 342536 236348
rect 342530 236308 342536 236320
rect 342588 236348 342594 236360
rect 416130 236348 416136 236360
rect 342588 236320 416136 236348
rect 342588 236308 342594 236320
rect 416130 236308 416136 236320
rect 416188 236308 416194 236360
rect 61372 236283 61430 236289
rect 61372 236249 61384 236283
rect 61418 236280 61430 236283
rect 61470 236280 61476 236292
rect 61418 236252 61476 236280
rect 61418 236249 61430 236252
rect 61372 236243 61430 236249
rect 61470 236240 61476 236252
rect 61528 236240 61534 236292
rect 342266 236283 342324 236289
rect 342266 236249 342278 236283
rect 342312 236249 342324 236283
rect 342266 236243 342324 236249
rect 62482 236212 62488 236224
rect 62443 236184 62488 236212
rect 62482 236172 62488 236184
rect 62540 236212 62546 236224
rect 155954 236212 155960 236224
rect 62540 236184 155960 236212
rect 62540 236172 62546 236184
rect 155954 236172 155960 236184
rect 156012 236172 156018 236224
rect 341150 236212 341156 236224
rect 341111 236184 341156 236212
rect 341150 236172 341156 236184
rect 341208 236172 341214 236224
rect 342272 236212 342300 236243
rect 342346 236212 342352 236224
rect 342272 236184 342352 236212
rect 342346 236172 342352 236184
rect 342404 236172 342410 236224
rect 240318 232472 240324 232484
rect 240279 232444 240324 232472
rect 240318 232432 240324 232444
rect 240376 232432 240382 232484
rect 216214 231520 216220 231532
rect 216175 231492 216220 231520
rect 216214 231480 216220 231492
rect 216272 231480 216278 231532
rect 418525 231047 418583 231053
rect 418525 231044 418537 231047
rect 412606 231016 418537 231044
rect 204346 230800 204352 230852
rect 204404 230840 204410 230852
rect 412606 230840 412634 231016
rect 418525 231013 418537 231016
rect 418571 231013 418583 231047
rect 418525 231007 418583 231013
rect 419074 230976 419080 230988
rect 419035 230948 419080 230976
rect 419074 230936 419080 230948
rect 419132 230976 419138 230988
rect 444190 230976 444196 230988
rect 419132 230948 444196 230976
rect 419132 230936 419138 230948
rect 444190 230936 444196 230948
rect 444248 230936 444254 230988
rect 418893 230843 418951 230849
rect 418893 230840 418905 230843
rect 204404 230812 412634 230840
rect 413112 230812 418905 230840
rect 204404 230800 204410 230812
rect 126974 230732 126980 230784
rect 127032 230772 127038 230784
rect 413112 230772 413140 230812
rect 418893 230809 418905 230812
rect 418939 230809 418951 230843
rect 418893 230803 418951 230809
rect 127032 230744 413140 230772
rect 127032 230732 127038 230744
rect 418706 230732 418712 230784
rect 418764 230772 418770 230784
rect 418985 230775 419043 230781
rect 418985 230772 418997 230775
rect 418764 230744 418997 230772
rect 418764 230732 418770 230744
rect 418985 230741 418997 230744
rect 419031 230741 419043 230775
rect 418985 230735 419043 230741
rect 153378 229820 153384 229832
rect 153339 229792 153384 229820
rect 153378 229780 153384 229792
rect 153436 229780 153442 229832
rect 153470 229780 153476 229832
rect 153528 229820 153534 229832
rect 153528 229792 153573 229820
rect 153528 229780 153534 229792
rect 167822 228392 167828 228404
rect 167783 228364 167828 228392
rect 167822 228352 167828 228364
rect 167880 228352 167886 228404
rect 167454 228256 167460 228268
rect 167415 228228 167460 228256
rect 167454 228216 167460 228228
rect 167512 228216 167518 228268
rect 167178 228188 167184 228200
rect 167139 228160 167184 228188
rect 167178 228148 167184 228160
rect 167236 228148 167242 228200
rect 167362 228188 167368 228200
rect 167323 228160 167368 228188
rect 167362 228148 167368 228160
rect 167420 228148 167426 228200
rect 175826 228188 175832 228200
rect 171106 228160 175832 228188
rect 167196 228120 167224 228148
rect 171106 228120 171134 228160
rect 175826 228148 175832 228160
rect 175884 228188 175890 228200
rect 180794 228188 180800 228200
rect 175884 228160 180800 228188
rect 175884 228148 175890 228160
rect 180794 228148 180800 228160
rect 180852 228148 180858 228200
rect 167196 228092 171134 228120
rect 292209 228055 292267 228061
rect 292209 228021 292221 228055
rect 292255 228052 292267 228055
rect 315574 228052 315580 228064
rect 292255 228024 315580 228052
rect 292255 228021 292267 228024
rect 292209 228015 292267 228021
rect 315574 228012 315580 228024
rect 315632 228012 315638 228064
rect 137186 227712 137192 227724
rect 137147 227684 137192 227712
rect 137186 227672 137192 227684
rect 137244 227672 137250 227724
rect 167638 227672 167644 227724
rect 167696 227712 167702 227724
rect 329742 227712 329748 227724
rect 167696 227684 329748 227712
rect 167696 227672 167702 227684
rect 329742 227672 329748 227684
rect 329800 227672 329806 227724
rect 136453 227647 136511 227653
rect 136453 227613 136465 227647
rect 136499 227613 136511 227647
rect 136453 227607 136511 227613
rect 136468 227576 136496 227607
rect 137186 227576 137192 227588
rect 136468 227548 137192 227576
rect 137186 227536 137192 227548
rect 137244 227536 137250 227588
rect 136729 227307 136787 227313
rect 136729 227273 136741 227307
rect 136775 227273 136787 227307
rect 136729 227267 136787 227273
rect 135622 227168 135628 227180
rect 135583 227140 135628 227168
rect 135622 227128 135628 227140
rect 135680 227128 135686 227180
rect 135898 227168 135904 227180
rect 135859 227140 135904 227168
rect 135898 227128 135904 227140
rect 135956 227128 135962 227180
rect 135990 227128 135996 227180
rect 136048 227168 136054 227180
rect 136177 227171 136235 227177
rect 136048 227140 136093 227168
rect 136048 227128 136054 227140
rect 136177 227137 136189 227171
rect 136223 227168 136235 227171
rect 136744 227168 136772 227267
rect 175642 227236 175648 227248
rect 136223 227140 136772 227168
rect 137020 227208 175648 227236
rect 136223 227137 136235 227140
rect 136177 227131 136235 227137
rect 135809 227103 135867 227109
rect 135809 227069 135821 227103
rect 135855 227069 135867 227103
rect 135809 227063 135867 227069
rect 135824 227032 135852 227063
rect 136542 227060 136548 227112
rect 136600 227100 136606 227112
rect 137020 227100 137048 227208
rect 175642 227196 175648 227208
rect 175700 227196 175706 227248
rect 137186 227100 137192 227112
rect 136600 227072 137048 227100
rect 137147 227072 137192 227100
rect 136600 227060 136606 227072
rect 137186 227060 137192 227072
rect 137244 227060 137250 227112
rect 167638 227100 167644 227112
rect 142126 227072 167644 227100
rect 142126 227032 142154 227072
rect 167638 227060 167644 227072
rect 167696 227060 167702 227112
rect 135824 227004 142154 227032
rect 40586 226924 40592 226976
rect 40644 226964 40650 226976
rect 135533 226967 135591 226973
rect 135533 226964 135545 226967
rect 40644 226936 135545 226964
rect 40644 226924 40650 226936
rect 135533 226933 135545 226936
rect 135579 226933 135591 226967
rect 135533 226927 135591 226933
rect 347038 225672 347044 225684
rect 346999 225644 347044 225672
rect 347038 225632 347044 225644
rect 347096 225632 347102 225684
rect 290274 224992 290280 225004
rect 290187 224964 290280 224992
rect 290274 224952 290280 224964
rect 290332 224992 290338 225004
rect 335906 224992 335912 225004
rect 290332 224964 335912 224992
rect 290332 224952 290338 224964
rect 335906 224952 335912 224964
rect 335964 224952 335970 225004
rect 289814 224788 289820 224800
rect 289775 224760 289820 224788
rect 289814 224748 289820 224760
rect 289872 224748 289878 224800
rect 100846 224584 100852 224596
rect 100807 224556 100852 224584
rect 100846 224544 100852 224556
rect 100904 224544 100910 224596
rect 289998 224584 290004 224596
rect 289959 224556 290004 224584
rect 289998 224544 290004 224556
rect 290056 224544 290062 224596
rect 289449 224451 289507 224457
rect 289449 224417 289461 224451
rect 289495 224448 289507 224451
rect 289814 224448 289820 224460
rect 289495 224420 289820 224448
rect 289495 224417 289507 224420
rect 289449 224411 289507 224417
rect 289814 224408 289820 224420
rect 289872 224408 289878 224460
rect 100938 224380 100944 224392
rect 100851 224352 100944 224380
rect 100938 224340 100944 224352
rect 100996 224380 101002 224392
rect 310790 224380 310796 224392
rect 100996 224352 310796 224380
rect 100996 224340 101002 224352
rect 310790 224340 310796 224352
rect 310848 224340 310854 224392
rect 32766 224204 32772 224256
rect 32824 224244 32830 224256
rect 289541 224247 289599 224253
rect 289541 224244 289553 224247
rect 32824 224216 289553 224244
rect 32824 224204 32830 224216
rect 289541 224213 289553 224216
rect 289587 224213 289599 224247
rect 289541 224207 289599 224213
rect 289630 224204 289636 224256
rect 289688 224244 289694 224256
rect 289688 224216 289733 224244
rect 289688 224204 289694 224216
rect 3050 223728 3056 223780
rect 3108 223768 3114 223780
rect 5902 223768 5908 223780
rect 3108 223740 5908 223768
rect 3108 223728 3114 223740
rect 5902 223728 5908 223740
rect 5960 223728 5966 223780
rect 227640 223672 228220 223700
rect 126974 223524 126980 223576
rect 127032 223564 127038 223576
rect 127526 223564 127532 223576
rect 127032 223536 127532 223564
rect 127032 223524 127038 223536
rect 127526 223524 127532 223536
rect 127584 223524 127590 223576
rect 141418 223524 141424 223576
rect 141476 223564 141482 223576
rect 142062 223564 142068 223576
rect 141476 223536 142068 223564
rect 141476 223524 141482 223536
rect 142062 223524 142068 223536
rect 142120 223524 142126 223576
rect 134518 223456 134524 223508
rect 134576 223496 134582 223508
rect 227640 223496 227668 223672
rect 228082 223564 228088 223576
rect 228008 223536 228088 223564
rect 134576 223468 227668 223496
rect 227901 223499 227959 223505
rect 134576 223456 134582 223468
rect 227901 223465 227913 223499
rect 227947 223496 227959 223499
rect 228008 223496 228036 223536
rect 228082 223524 228088 223536
rect 228140 223524 228146 223576
rect 227947 223468 228036 223496
rect 228192 223496 228220 223672
rect 260834 223524 260840 223576
rect 260892 223564 260898 223576
rect 265713 223567 265771 223573
rect 265713 223564 265725 223567
rect 260892 223536 265725 223564
rect 260892 223524 260898 223536
rect 265713 223533 265725 223536
rect 265759 223533 265771 223567
rect 265713 223527 265771 223533
rect 467650 223496 467656 223508
rect 228192 223468 467656 223496
rect 227947 223465 227959 223468
rect 227901 223459 227959 223465
rect 467650 223456 467656 223468
rect 467708 223456 467714 223508
rect 207382 223388 207388 223440
rect 207440 223428 207446 223440
rect 379514 223428 379520 223440
rect 207440 223400 379520 223428
rect 207440 223388 207446 223400
rect 379514 223388 379520 223400
rect 379572 223388 379578 223440
rect 42058 223320 42064 223372
rect 42116 223360 42122 223372
rect 239030 223360 239036 223372
rect 42116 223332 239036 223360
rect 42116 223320 42122 223332
rect 239030 223320 239036 223332
rect 239088 223320 239094 223372
rect 265713 223363 265771 223369
rect 248386 223332 263594 223360
rect 187602 223252 187608 223304
rect 187660 223292 187666 223304
rect 248386 223292 248414 223332
rect 260466 223292 260472 223304
rect 187660 223264 248414 223292
rect 260427 223264 260472 223292
rect 187660 223252 187666 223264
rect 260466 223252 260472 223264
rect 260524 223252 260530 223304
rect 260558 223252 260564 223304
rect 260616 223292 260622 223304
rect 260837 223295 260895 223301
rect 260837 223292 260849 223295
rect 260616 223264 260849 223292
rect 260616 223252 260622 223264
rect 260837 223261 260849 223264
rect 260883 223261 260895 223295
rect 263566 223292 263594 223332
rect 265713 223329 265725 223363
rect 265759 223360 265771 223363
rect 367278 223360 367284 223372
rect 265759 223332 367284 223360
rect 265759 223329 265771 223332
rect 265713 223323 265771 223329
rect 367278 223320 367284 223332
rect 367336 223320 367342 223372
rect 430574 223292 430580 223304
rect 263566 223264 430580 223292
rect 260837 223255 260895 223261
rect 430574 223252 430580 223264
rect 430632 223252 430638 223304
rect 194410 223184 194416 223236
rect 194468 223224 194474 223236
rect 255958 223224 255964 223236
rect 194468 223196 255964 223224
rect 194468 223184 194474 223196
rect 255958 223184 255964 223196
rect 256016 223184 256022 223236
rect 260742 223184 260748 223236
rect 260800 223224 260806 223236
rect 496630 223224 496636 223236
rect 260800 223196 496636 223224
rect 260800 223184 260806 223196
rect 496630 223184 496636 223196
rect 496688 223184 496694 223236
rect 61838 223116 61844 223168
rect 61896 223156 61902 223168
rect 260558 223156 260564 223168
rect 61896 223128 260564 223156
rect 61896 223116 61902 223128
rect 260558 223116 260564 223128
rect 260616 223116 260622 223168
rect 260650 223116 260656 223168
rect 260708 223156 260714 223168
rect 260837 223159 260895 223165
rect 260708 223128 260753 223156
rect 260708 223116 260714 223128
rect 260837 223125 260849 223159
rect 260883 223156 260895 223159
rect 382274 223156 382280 223168
rect 260883 223128 382280 223156
rect 260883 223125 260895 223128
rect 260837 223119 260895 223125
rect 382274 223116 382280 223128
rect 382332 223116 382338 223168
rect 93670 223048 93676 223100
rect 93728 223088 93734 223100
rect 147766 223088 147772 223100
rect 93728 223060 147772 223088
rect 93728 223048 93734 223060
rect 147766 223048 147772 223060
rect 147824 223048 147830 223100
rect 112254 222980 112260 223032
rect 112312 223020 112318 223032
rect 200390 223020 200396 223032
rect 112312 222992 200396 223020
rect 112312 222980 112318 222992
rect 200390 222980 200396 222992
rect 200448 222980 200454 223032
rect 280522 222980 280528 223032
rect 280580 223020 280586 223032
rect 328454 223020 328460 223032
rect 280580 222992 328460 223020
rect 280580 222980 280586 222992
rect 328454 222980 328460 222992
rect 328512 222980 328518 223032
rect 35158 222912 35164 222964
rect 35216 222952 35222 222964
rect 426802 222952 426808 222964
rect 35216 222924 426808 222952
rect 35216 222912 35222 222924
rect 426802 222912 426808 222924
rect 426860 222912 426866 222964
rect 95050 222844 95056 222896
rect 95108 222884 95114 222896
rect 496354 222884 496360 222896
rect 95108 222856 496360 222884
rect 95108 222844 95114 222856
rect 496354 222844 496360 222856
rect 496412 222844 496418 222896
rect 81802 222776 81808 222828
rect 81860 222816 81866 222828
rect 82722 222816 82728 222828
rect 81860 222788 82728 222816
rect 81860 222776 81866 222788
rect 82722 222776 82728 222788
rect 82780 222776 82786 222828
rect 140866 222776 140872 222828
rect 140924 222816 140930 222828
rect 247126 222816 247132 222828
rect 140924 222788 247132 222816
rect 140924 222776 140930 222788
rect 247126 222776 247132 222788
rect 247184 222776 247190 222828
rect 199930 222708 199936 222760
rect 199988 222748 199994 222760
rect 299750 222748 299756 222760
rect 199988 222720 299756 222748
rect 199988 222708 199994 222720
rect 299750 222708 299756 222720
rect 299808 222708 299814 222760
rect 53834 222640 53840 222692
rect 53892 222680 53898 222692
rect 54662 222680 54668 222692
rect 53892 222652 54668 222680
rect 53892 222640 53898 222652
rect 54662 222640 54668 222652
rect 54720 222640 54726 222692
rect 153194 222640 153200 222692
rect 153252 222680 153258 222692
rect 154022 222680 154028 222692
rect 153252 222652 154028 222680
rect 153252 222640 153258 222652
rect 154022 222640 154028 222652
rect 154080 222640 154086 222692
rect 205818 222640 205824 222692
rect 205876 222680 205882 222692
rect 286502 222680 286508 222692
rect 205876 222652 286508 222680
rect 205876 222640 205882 222652
rect 286502 222640 286508 222652
rect 286560 222640 286566 222692
rect 101398 222572 101404 222624
rect 101456 222612 101462 222624
rect 438486 222612 438492 222624
rect 101456 222584 438492 222612
rect 101456 222572 101462 222584
rect 438486 222572 438492 222584
rect 438544 222572 438550 222624
rect 252554 222504 252560 222556
rect 252612 222544 252618 222556
rect 253382 222544 253388 222556
rect 252612 222516 253388 222544
rect 252612 222504 252618 222516
rect 253382 222504 253388 222516
rect 253440 222504 253446 222556
rect 68554 222368 68560 222420
rect 68612 222408 68618 222420
rect 259178 222408 259184 222420
rect 68612 222380 259184 222408
rect 68612 222368 68618 222380
rect 259178 222368 259184 222380
rect 259236 222368 259242 222420
rect 260650 222368 260656 222420
rect 260708 222408 260714 222420
rect 475378 222408 475384 222420
rect 260708 222380 475384 222408
rect 260708 222368 260714 222380
rect 475378 222368 475384 222380
rect 475436 222368 475442 222420
rect 227530 222300 227536 222352
rect 227588 222340 227594 222352
rect 496722 222340 496728 222352
rect 227588 222312 496728 222340
rect 227588 222300 227594 222312
rect 496722 222300 496728 222312
rect 496780 222300 496786 222352
rect 7190 222232 7196 222284
rect 7248 222272 7254 222284
rect 21634 222272 21640 222284
rect 7248 222244 21640 222272
rect 7248 222232 7254 222244
rect 21634 222232 21640 222244
rect 21692 222232 21698 222284
rect 48682 222232 48688 222284
rect 48740 222272 48746 222284
rect 381078 222272 381084 222284
rect 48740 222244 381084 222272
rect 48740 222232 48746 222244
rect 381078 222232 381084 222244
rect 381136 222232 381142 222284
rect 15562 222164 15568 222216
rect 15620 222204 15626 222216
rect 362218 222204 362224 222216
rect 15620 222176 362224 222204
rect 15620 222164 15626 222176
rect 362218 222164 362224 222176
rect 362276 222164 362282 222216
rect 79778 220776 79784 220788
rect 79739 220748 79784 220776
rect 79778 220736 79784 220748
rect 79836 220736 79842 220788
rect 97074 220776 97080 220788
rect 97035 220748 97080 220776
rect 97074 220736 97080 220748
rect 97132 220736 97138 220788
rect 123386 220776 123392 220788
rect 123347 220748 123392 220776
rect 123386 220736 123392 220748
rect 123444 220736 123450 220788
rect 131853 220779 131911 220785
rect 131853 220745 131865 220779
rect 131899 220776 131911 220779
rect 164145 220779 164203 220785
rect 131899 220748 132494 220776
rect 131899 220745 131911 220748
rect 131853 220739 131911 220745
rect 112530 220708 112536 220720
rect 55186 220680 112536 220708
rect 50065 220643 50123 220649
rect 50065 220609 50077 220643
rect 50111 220640 50123 220643
rect 55186 220640 55214 220680
rect 112530 220668 112536 220680
rect 112588 220668 112594 220720
rect 128449 220711 128507 220717
rect 128449 220677 128461 220711
rect 128495 220708 128507 220711
rect 129645 220711 129703 220717
rect 129645 220708 129657 220711
rect 128495 220680 129657 220708
rect 128495 220677 128507 220680
rect 128449 220671 128507 220677
rect 129645 220677 129657 220680
rect 129691 220677 129703 220711
rect 132466 220708 132494 220748
rect 164145 220745 164157 220779
rect 164191 220776 164203 220779
rect 164191 220748 171134 220776
rect 164191 220745 164203 220748
rect 164145 220739 164203 220745
rect 159082 220708 159088 220720
rect 132466 220680 159088 220708
rect 129645 220671 129703 220677
rect 159082 220668 159088 220680
rect 159140 220668 159146 220720
rect 171106 220708 171134 220748
rect 204990 220736 204996 220788
rect 205048 220776 205054 220788
rect 205450 220776 205456 220788
rect 205048 220748 205456 220776
rect 205048 220736 205054 220748
rect 205450 220736 205456 220748
rect 205508 220736 205514 220788
rect 205634 220776 205640 220788
rect 205595 220748 205640 220776
rect 205634 220736 205640 220748
rect 205692 220736 205698 220788
rect 205726 220736 205732 220788
rect 205784 220776 205790 220788
rect 209038 220776 209044 220788
rect 205784 220748 209044 220776
rect 205784 220736 205790 220748
rect 209038 220736 209044 220748
rect 209096 220776 209102 220788
rect 341242 220776 341248 220788
rect 209096 220748 341248 220776
rect 209096 220736 209102 220748
rect 341242 220736 341248 220748
rect 341300 220736 341306 220788
rect 248690 220708 248696 220720
rect 171106 220680 248696 220708
rect 248690 220668 248696 220680
rect 248748 220708 248754 220720
rect 249702 220708 249708 220720
rect 248748 220680 249708 220708
rect 248748 220668 248754 220680
rect 249702 220668 249708 220680
rect 249760 220668 249766 220720
rect 258902 220708 258908 220720
rect 251376 220680 258908 220708
rect 50111 220612 55214 220640
rect 75733 220643 75791 220649
rect 50111 220609 50123 220612
rect 50065 220603 50123 220609
rect 75733 220609 75745 220643
rect 75779 220640 75791 220643
rect 75825 220643 75883 220649
rect 75825 220640 75837 220643
rect 75779 220612 75837 220640
rect 75779 220609 75791 220612
rect 75733 220603 75791 220609
rect 75825 220609 75837 220612
rect 75871 220609 75883 220643
rect 79410 220640 79416 220652
rect 79371 220612 79416 220640
rect 75825 220603 75883 220609
rect 79410 220600 79416 220612
rect 79468 220600 79474 220652
rect 96709 220643 96767 220649
rect 96709 220609 96721 220643
rect 96755 220640 96767 220643
rect 107654 220640 107660 220652
rect 96755 220612 107660 220640
rect 96755 220609 96767 220612
rect 96709 220603 96767 220609
rect 107654 220600 107660 220612
rect 107712 220600 107718 220652
rect 123481 220643 123539 220649
rect 123481 220609 123493 220643
rect 123527 220640 123539 220643
rect 124125 220643 124183 220649
rect 124125 220640 124137 220643
rect 123527 220612 124137 220640
rect 123527 220609 123539 220612
rect 123481 220603 123539 220609
rect 124125 220609 124137 220612
rect 124171 220609 124183 220643
rect 124125 220603 124183 220609
rect 128357 220643 128415 220649
rect 128357 220609 128369 220643
rect 128403 220640 128415 220643
rect 129553 220643 129611 220649
rect 129553 220640 129565 220643
rect 128403 220612 129565 220640
rect 128403 220609 128415 220612
rect 128357 220603 128415 220609
rect 129553 220609 129565 220612
rect 129599 220609 129611 220643
rect 129553 220603 129611 220609
rect 132977 220643 133035 220649
rect 132977 220609 132989 220643
rect 133023 220640 133035 220643
rect 133785 220643 133843 220649
rect 133785 220640 133797 220643
rect 133023 220612 133797 220640
rect 133023 220609 133035 220612
rect 132977 220603 133035 220609
rect 133785 220609 133797 220612
rect 133831 220609 133843 220643
rect 133785 220603 133843 220609
rect 163032 220643 163090 220649
rect 163032 220609 163044 220643
rect 163078 220640 163090 220643
rect 167089 220643 167147 220649
rect 167089 220640 167101 220643
rect 163078 220612 167101 220640
rect 163078 220609 163090 220612
rect 163032 220603 163090 220609
rect 167089 220609 167101 220612
rect 167135 220609 167147 220643
rect 178310 220640 178316 220652
rect 178271 220612 178316 220640
rect 167089 220603 167147 220609
rect 178310 220600 178316 220612
rect 178368 220600 178374 220652
rect 204990 220640 204996 220652
rect 204951 220612 204996 220640
rect 204990 220600 204996 220612
rect 205048 220600 205054 220652
rect 205174 220640 205180 220652
rect 205135 220612 205180 220640
rect 205174 220600 205180 220612
rect 205232 220600 205238 220652
rect 205266 220600 205272 220652
rect 205324 220640 205330 220652
rect 205545 220643 205603 220649
rect 205545 220640 205557 220643
rect 205324 220612 205369 220640
rect 205468 220612 205557 220640
rect 205324 220600 205330 220612
rect 78953 220575 79011 220581
rect 78953 220541 78965 220575
rect 78999 220572 79011 220575
rect 79137 220575 79195 220581
rect 79137 220572 79149 220575
rect 78999 220544 79149 220572
rect 78999 220541 79011 220544
rect 78953 220535 79011 220541
rect 79137 220541 79149 220544
rect 79183 220541 79195 220575
rect 79318 220572 79324 220584
rect 79279 220544 79324 220572
rect 79137 220535 79195 220541
rect 79318 220532 79324 220544
rect 79376 220532 79382 220584
rect 96157 220575 96215 220581
rect 96157 220541 96169 220575
rect 96203 220572 96215 220575
rect 96433 220575 96491 220581
rect 96433 220572 96445 220575
rect 96203 220544 96445 220572
rect 96203 220541 96215 220544
rect 96157 220535 96215 220541
rect 96433 220541 96445 220544
rect 96479 220541 96491 220575
rect 96614 220572 96620 220584
rect 96575 220544 96620 220572
rect 96433 220535 96491 220541
rect 96614 220532 96620 220544
rect 96672 220532 96678 220584
rect 97169 220575 97227 220581
rect 97169 220541 97181 220575
rect 97215 220572 97227 220575
rect 129093 220575 129151 220581
rect 129093 220572 129105 220575
rect 97215 220544 129105 220572
rect 97215 220541 97227 220544
rect 97169 220535 97227 220541
rect 129093 220541 129105 220544
rect 129139 220572 129151 220575
rect 129369 220575 129427 220581
rect 129369 220572 129381 220575
rect 129139 220544 129381 220572
rect 129139 220541 129151 220544
rect 129093 220535 129151 220541
rect 129369 220541 129381 220544
rect 129415 220541 129427 220575
rect 129369 220535 129427 220541
rect 133230 220532 133236 220584
rect 133288 220572 133294 220584
rect 162762 220572 162768 220584
rect 133288 220544 133381 220572
rect 142126 220544 162768 220572
rect 133288 220532 133294 220544
rect 55030 220504 55036 220516
rect 54991 220476 55036 220504
rect 55030 220464 55036 220476
rect 55088 220464 55094 220516
rect 75641 220507 75699 220513
rect 75641 220473 75653 220507
rect 75687 220504 75699 220507
rect 125778 220504 125784 220516
rect 75687 220476 125784 220504
rect 75687 220473 75699 220476
rect 75641 220467 75699 220473
rect 125778 220464 125784 220476
rect 125836 220464 125842 220516
rect 133248 220504 133276 220532
rect 137922 220504 137928 220516
rect 133248 220476 137928 220504
rect 137922 220464 137928 220476
rect 137980 220504 137986 220516
rect 142126 220504 142154 220544
rect 162762 220532 162768 220544
rect 162820 220532 162826 220584
rect 205358 220572 205364 220584
rect 205319 220544 205364 220572
rect 205358 220532 205364 220544
rect 205416 220532 205422 220584
rect 205468 220572 205496 220612
rect 205545 220609 205557 220612
rect 205591 220609 205603 220643
rect 235258 220640 235264 220652
rect 235219 220612 235264 220640
rect 205545 220603 205603 220609
rect 235258 220600 235264 220612
rect 235316 220600 235322 220652
rect 251376 220572 251404 220680
rect 258902 220668 258908 220680
rect 258960 220668 258966 220720
rect 259270 220708 259276 220720
rect 259231 220680 259276 220708
rect 259270 220668 259276 220680
rect 259328 220668 259334 220720
rect 266078 220668 266084 220720
rect 266136 220668 266142 220720
rect 266633 220711 266691 220717
rect 266633 220677 266645 220711
rect 266679 220708 266691 220711
rect 430942 220708 430948 220720
rect 266679 220680 430948 220708
rect 266679 220677 266691 220680
rect 266633 220671 266691 220677
rect 430942 220668 430948 220680
rect 431000 220668 431006 220720
rect 257430 220640 257436 220652
rect 257391 220612 257436 220640
rect 257430 220600 257436 220612
rect 257488 220600 257494 220652
rect 259086 220649 259092 220652
rect 257525 220643 257583 220649
rect 257525 220609 257537 220643
rect 257571 220640 257583 220643
rect 257985 220643 258043 220649
rect 257985 220640 257997 220643
rect 257571 220612 257997 220640
rect 257571 220609 257583 220612
rect 257525 220603 257583 220609
rect 257985 220609 257997 220612
rect 258031 220609 258043 220643
rect 259084 220640 259092 220649
rect 259047 220612 259092 220640
rect 257985 220603 258043 220609
rect 259084 220603 259092 220612
rect 259086 220600 259092 220603
rect 259144 220600 259150 220652
rect 259178 220600 259184 220652
rect 259236 220640 259242 220652
rect 259454 220640 259460 220652
rect 259236 220612 259281 220640
rect 259415 220612 259460 220640
rect 259236 220600 259242 220612
rect 259454 220600 259460 220612
rect 259512 220600 259518 220652
rect 259549 220643 259607 220649
rect 259549 220609 259561 220643
rect 259595 220640 259607 220643
rect 259638 220640 259644 220652
rect 259595 220612 259644 220640
rect 259595 220609 259607 220612
rect 259549 220603 259607 220609
rect 259638 220600 259644 220612
rect 259696 220600 259702 220652
rect 266096 220640 266124 220668
rect 263566 220612 266124 220640
rect 266193 220643 266251 220649
rect 257154 220572 257160 220584
rect 205468 220544 251404 220572
rect 257115 220544 257160 220572
rect 137980 220476 142154 220504
rect 204809 220507 204867 220513
rect 137980 220464 137986 220476
rect 204809 220473 204821 220507
rect 204855 220504 204867 220507
rect 205468 220504 205496 220544
rect 257154 220532 257160 220544
rect 257212 220532 257218 220584
rect 257246 220532 257252 220584
rect 257304 220572 257310 220584
rect 263566 220572 263594 220612
rect 266193 220609 266205 220643
rect 266239 220640 266251 220643
rect 267001 220643 267059 220649
rect 266239 220612 266952 220640
rect 266239 220609 266251 220612
rect 266193 220603 266251 220609
rect 257304 220544 257349 220572
rect 257540 220544 263594 220572
rect 266449 220575 266507 220581
rect 257304 220532 257310 220544
rect 204855 220476 205496 220504
rect 204855 220473 204867 220476
rect 204809 220467 204867 220473
rect 205542 220464 205548 220516
rect 205600 220504 205606 220516
rect 257338 220504 257344 220516
rect 205600 220476 257344 220504
rect 205600 220464 205606 220476
rect 257338 220464 257344 220476
rect 257396 220464 257402 220516
rect 49970 220436 49976 220448
rect 49931 220408 49976 220436
rect 49970 220396 49976 220408
rect 50028 220396 50034 220448
rect 75825 220439 75883 220445
rect 75825 220405 75837 220439
rect 75871 220405 75883 220439
rect 77754 220436 77760 220448
rect 77715 220408 77760 220436
rect 75825 220399 75883 220405
rect 75840 220232 75868 220399
rect 77754 220396 77760 220408
rect 77812 220396 77818 220448
rect 78953 220439 79011 220445
rect 78953 220405 78965 220439
rect 78999 220436 79011 220439
rect 96157 220439 96215 220445
rect 96157 220436 96169 220439
rect 78999 220408 96169 220436
rect 78999 220405 79011 220408
rect 78953 220399 79011 220405
rect 96157 220405 96169 220408
rect 96203 220436 96215 220439
rect 97169 220439 97227 220445
rect 97169 220436 97181 220439
rect 96203 220408 97181 220436
rect 96203 220405 96215 220408
rect 96157 220399 96215 220405
rect 97169 220405 97181 220408
rect 97215 220405 97227 220439
rect 97169 220399 97227 220405
rect 130013 220439 130071 220445
rect 130013 220405 130025 220439
rect 130059 220436 130071 220439
rect 178037 220439 178095 220445
rect 130059 220408 131252 220436
rect 130059 220405 130071 220408
rect 130013 220399 130071 220405
rect 125318 220232 125324 220244
rect 75840 220204 125324 220232
rect 125318 220192 125324 220204
rect 125376 220192 125382 220244
rect 131224 220232 131252 220408
rect 178037 220405 178049 220439
rect 178083 220436 178095 220439
rect 178405 220439 178463 220445
rect 178405 220436 178417 220439
rect 178083 220408 178417 220436
rect 178083 220405 178095 220408
rect 178037 220399 178095 220405
rect 178405 220405 178417 220408
rect 178451 220405 178463 220439
rect 178405 220399 178463 220405
rect 205266 220396 205272 220448
rect 205324 220436 205330 220448
rect 213178 220436 213184 220448
rect 205324 220408 213184 220436
rect 205324 220396 205330 220408
rect 213178 220396 213184 220408
rect 213236 220436 213242 220448
rect 257540 220436 257568 220544
rect 266449 220541 266461 220575
rect 266495 220572 266507 220575
rect 266630 220572 266636 220584
rect 266495 220544 266636 220572
rect 266495 220541 266507 220544
rect 266449 220535 266507 220541
rect 266630 220532 266636 220544
rect 266688 220532 266694 220584
rect 266924 220572 266952 220612
rect 267001 220609 267013 220643
rect 267047 220640 267059 220643
rect 282914 220640 282920 220652
rect 267047 220612 282920 220640
rect 267047 220609 267059 220612
rect 267001 220603 267059 220609
rect 282914 220600 282920 220612
rect 282972 220600 282978 220652
rect 287609 220643 287667 220649
rect 287609 220609 287621 220643
rect 287655 220640 287667 220643
rect 288253 220643 288311 220649
rect 288253 220640 288265 220643
rect 287655 220612 288265 220640
rect 287655 220609 287667 220612
rect 287609 220603 287667 220609
rect 288253 220609 288265 220612
rect 288299 220609 288311 220643
rect 288253 220603 288311 220609
rect 272429 220575 272487 220581
rect 272429 220572 272441 220575
rect 266924 220544 272441 220572
rect 272429 220541 272441 220544
rect 272475 220541 272487 220575
rect 272429 220535 272487 220541
rect 272521 220575 272579 220581
rect 272521 220541 272533 220575
rect 272567 220572 272579 220575
rect 342530 220572 342536 220584
rect 272567 220544 342536 220572
rect 272567 220541 272579 220544
rect 272521 220535 272579 220541
rect 342530 220532 342536 220544
rect 342588 220532 342594 220584
rect 257614 220464 257620 220516
rect 257672 220504 257678 220516
rect 318518 220504 318524 220516
rect 257672 220476 265204 220504
rect 257672 220464 257678 220476
rect 257706 220436 257712 220448
rect 213236 220408 257568 220436
rect 257667 220408 257712 220436
rect 213236 220396 213242 220408
rect 257706 220396 257712 220408
rect 257764 220396 257770 220448
rect 258077 220439 258135 220445
rect 258077 220405 258089 220439
rect 258123 220436 258135 220439
rect 258905 220439 258963 220445
rect 258905 220436 258917 220439
rect 258123 220408 258917 220436
rect 258123 220405 258135 220408
rect 258077 220399 258135 220405
rect 258905 220405 258917 220408
rect 258951 220405 258963 220439
rect 265066 220436 265072 220448
rect 265027 220408 265072 220436
rect 258905 220399 258963 220405
rect 265066 220396 265072 220408
rect 265124 220396 265130 220448
rect 265176 220436 265204 220476
rect 266464 220476 318524 220504
rect 266464 220436 266492 220476
rect 318518 220464 318524 220476
rect 318576 220464 318582 220516
rect 265176 220408 266492 220436
rect 266538 220396 266544 220448
rect 266596 220436 266602 220448
rect 341334 220436 341340 220448
rect 266596 220408 341340 220436
rect 266596 220396 266602 220408
rect 341334 220396 341340 220408
rect 341392 220396 341398 220448
rect 266630 220328 266636 220380
rect 266688 220368 266694 220380
rect 272521 220371 272579 220377
rect 272521 220368 272533 220371
rect 266688 220340 272533 220368
rect 266688 220328 266694 220340
rect 272521 220337 272533 220340
rect 272567 220337 272579 220371
rect 272521 220331 272579 220337
rect 317230 220232 317236 220244
rect 131224 220204 317236 220232
rect 317230 220192 317236 220204
rect 317288 220192 317294 220244
rect 133785 220167 133843 220173
rect 133785 220133 133797 220167
rect 133831 220164 133843 220167
rect 315666 220164 315672 220176
rect 133831 220136 315672 220164
rect 133831 220133 133843 220136
rect 133785 220127 133843 220133
rect 315666 220124 315672 220136
rect 315724 220124 315730 220176
rect 318702 220124 318708 220176
rect 318760 220164 318766 220176
rect 361666 220164 361672 220176
rect 318760 220136 361672 220164
rect 318760 220124 318766 220136
rect 361666 220124 361672 220136
rect 361724 220124 361730 220176
rect 23014 220056 23020 220108
rect 23072 220096 23078 220108
rect 178037 220099 178095 220105
rect 178037 220096 178049 220099
rect 23072 220068 178049 220096
rect 23072 220056 23078 220068
rect 178037 220065 178049 220068
rect 178083 220065 178095 220099
rect 178037 220059 178095 220065
rect 238478 220056 238484 220108
rect 238536 220096 238542 220108
rect 258077 220099 258135 220105
rect 258077 220096 258089 220099
rect 238536 220068 258089 220096
rect 238536 220056 238542 220068
rect 258077 220065 258089 220068
rect 258123 220065 258135 220099
rect 258077 220059 258135 220065
rect 259638 220056 259644 220108
rect 259696 220096 259702 220108
rect 267001 220099 267059 220105
rect 267001 220096 267013 220099
rect 259696 220068 267013 220096
rect 259696 220056 259702 220068
rect 267001 220065 267013 220068
rect 267047 220065 267059 220099
rect 267001 220059 267059 220065
rect 272429 220099 272487 220105
rect 272429 220065 272441 220099
rect 272475 220096 272487 220099
rect 340414 220096 340420 220108
rect 272475 220068 340420 220096
rect 272475 220065 272487 220068
rect 272429 220059 272487 220065
rect 340414 220056 340420 220068
rect 340472 220056 340478 220108
rect 167089 220031 167147 220037
rect 167089 219997 167101 220031
rect 167135 220028 167147 220031
rect 310606 220028 310612 220040
rect 167135 220000 310612 220028
rect 167135 219997 167147 220000
rect 167089 219991 167147 219997
rect 310606 219988 310612 220000
rect 310664 219988 310670 220040
rect 129093 219963 129151 219969
rect 129093 219929 129105 219963
rect 129139 219960 129151 219963
rect 167178 219960 167184 219972
rect 129139 219932 167184 219960
rect 129139 219929 129151 219932
rect 129093 219923 129151 219929
rect 167178 219920 167184 219932
rect 167236 219920 167242 219972
rect 257985 219963 258043 219969
rect 257985 219929 257997 219963
rect 258031 219960 258043 219963
rect 318334 219960 318340 219972
rect 258031 219932 318340 219960
rect 258031 219929 258043 219932
rect 257985 219923 258043 219929
rect 318334 219920 318340 219932
rect 318392 219920 318398 219972
rect 124125 219895 124183 219901
rect 124125 219861 124137 219895
rect 124171 219892 124183 219895
rect 204809 219895 204867 219901
rect 204809 219892 204821 219895
rect 124171 219864 204821 219892
rect 124171 219861 124183 219864
rect 124125 219855 124183 219861
rect 204809 219861 204821 219864
rect 204855 219861 204867 219895
rect 204809 219855 204867 219861
rect 259454 219852 259460 219904
rect 259512 219892 259518 219904
rect 266633 219895 266691 219901
rect 266633 219892 266645 219895
rect 259512 219864 266645 219892
rect 259512 219852 259518 219864
rect 266633 219861 266645 219864
rect 266679 219861 266691 219895
rect 266633 219855 266691 219861
rect 266725 219895 266783 219901
rect 266725 219861 266737 219895
rect 266771 219892 266783 219895
rect 318702 219892 318708 219904
rect 266771 219864 318708 219892
rect 266771 219861 266783 219864
rect 266725 219855 266783 219861
rect 318702 219852 318708 219864
rect 318760 219852 318766 219904
rect 254949 219827 255007 219833
rect 254949 219793 254961 219827
rect 254995 219824 255007 219827
rect 264974 219824 264980 219836
rect 254995 219796 264980 219824
rect 254995 219793 255007 219796
rect 254949 219787 255007 219793
rect 264974 219784 264980 219796
rect 265032 219784 265038 219836
rect 265066 219784 265072 219836
rect 265124 219824 265130 219836
rect 313182 219824 313188 219836
rect 265124 219796 313188 219824
rect 265124 219784 265130 219796
rect 313182 219784 313188 219796
rect 313240 219784 313246 219836
rect 249702 219716 249708 219768
rect 249760 219756 249766 219768
rect 310330 219756 310336 219768
rect 249760 219728 310336 219756
rect 249760 219716 249766 219728
rect 310330 219716 310336 219728
rect 310388 219716 310394 219768
rect 162762 219648 162768 219700
rect 162820 219688 162826 219700
rect 254949 219691 255007 219697
rect 254949 219688 254961 219691
rect 162820 219660 254961 219688
rect 162820 219648 162826 219660
rect 254949 219657 254961 219660
rect 254995 219657 255007 219691
rect 254949 219651 255007 219657
rect 259086 219648 259092 219700
rect 259144 219688 259150 219700
rect 266725 219691 266783 219697
rect 266725 219688 266737 219691
rect 259144 219660 266737 219688
rect 259144 219648 259150 219660
rect 266725 219657 266737 219660
rect 266771 219657 266783 219691
rect 266725 219651 266783 219657
rect 282914 219648 282920 219700
rect 282972 219688 282978 219700
rect 317138 219688 317144 219700
rect 282972 219660 317144 219688
rect 282972 219648 282978 219660
rect 317138 219648 317144 219660
rect 317196 219648 317202 219700
rect 205174 219580 205180 219632
rect 205232 219620 205238 219632
rect 495986 219620 495992 219632
rect 205232 219592 495992 219620
rect 205232 219580 205238 219592
rect 495986 219580 495992 219592
rect 496044 219580 496050 219632
rect 11790 219552 11796 219564
rect 11751 219524 11796 219552
rect 11790 219512 11796 219524
rect 11848 219512 11854 219564
rect 12802 219552 12808 219564
rect 12763 219524 12808 219552
rect 12802 219512 12808 219524
rect 12860 219512 12866 219564
rect 16206 219552 16212 219564
rect 16167 219524 16212 219552
rect 16206 219512 16212 219524
rect 16264 219512 16270 219564
rect 17218 219552 17224 219564
rect 17179 219524 17224 219552
rect 17218 219512 17224 219524
rect 17276 219512 17282 219564
rect 96062 219552 96068 219564
rect 45526 219524 55214 219552
rect 96023 219524 96068 219552
rect 4430 219444 4436 219496
rect 4488 219484 4494 219496
rect 45526 219484 45554 219524
rect 53742 219484 53748 219496
rect 4488 219456 45554 219484
rect 53703 219456 53748 219484
rect 4488 219444 4494 219456
rect 53742 219444 53748 219456
rect 53800 219444 53806 219496
rect 55186 219484 55214 219524
rect 96062 219512 96068 219524
rect 96120 219512 96126 219564
rect 257154 219512 257160 219564
rect 257212 219552 257218 219564
rect 318426 219552 318432 219564
rect 257212 219524 318432 219552
rect 257212 219512 257218 219524
rect 318426 219512 318432 219524
rect 318484 219512 318490 219564
rect 287609 219487 287667 219493
rect 287609 219484 287621 219487
rect 55186 219456 287621 219484
rect 287609 219453 287621 219456
rect 287655 219453 287667 219487
rect 287609 219447 287667 219453
rect 3602 219376 3608 219428
rect 3660 219416 3666 219428
rect 130378 219416 130384 219428
rect 3660 219388 130384 219416
rect 3660 219376 3666 219388
rect 130378 219376 130384 219388
rect 130436 219376 130442 219428
rect 7834 219308 7840 219360
rect 7892 219348 7898 219360
rect 20530 219348 20536 219360
rect 7892 219320 20536 219348
rect 7892 219308 7898 219320
rect 20530 219308 20536 219320
rect 20588 219308 20594 219360
rect 21542 219308 21548 219360
rect 21600 219308 21606 219360
rect 22922 219348 22928 219360
rect 22883 219320 22928 219348
rect 22922 219308 22928 219320
rect 22980 219308 22986 219360
rect 55490 219348 55496 219360
rect 45526 219320 55496 219348
rect 7742 219240 7748 219292
rect 7800 219280 7806 219292
rect 21560 219280 21588 219308
rect 7800 219252 21588 219280
rect 7800 219240 7806 219252
rect 8478 219172 8484 219224
rect 8536 219212 8542 219224
rect 45526 219212 45554 219320
rect 55490 219308 55496 219320
rect 55548 219308 55554 219360
rect 78122 219348 78128 219360
rect 78083 219320 78128 219348
rect 78122 219308 78128 219320
rect 78180 219308 78186 219360
rect 101490 219348 101496 219360
rect 84166 219320 101496 219348
rect 8536 219184 45554 219212
rect 8536 219172 8542 219184
rect 8202 219104 8208 219156
rect 8260 219144 8266 219156
rect 84166 219144 84194 219320
rect 101490 219308 101496 219320
rect 101548 219308 101554 219360
rect 112990 219348 112996 219360
rect 109006 219320 112996 219348
rect 8260 219116 84194 219144
rect 8260 219104 8266 219116
rect 9493 219079 9551 219085
rect 9493 219045 9505 219079
rect 9539 219076 9551 219079
rect 109006 219076 109034 219320
rect 112990 219308 112996 219320
rect 113048 219308 113054 219360
rect 114370 219348 114376 219360
rect 114331 219320 114376 219348
rect 114370 219308 114376 219320
rect 114428 219308 114434 219360
rect 218514 219308 218520 219360
rect 218572 219348 218578 219360
rect 232958 219348 232964 219360
rect 218572 219320 224954 219348
rect 232919 219320 232964 219348
rect 218572 219308 218578 219320
rect 9539 219048 109034 219076
rect 9539 219045 9551 219048
rect 9493 219039 9551 219045
rect 5442 218968 5448 219020
rect 5500 219008 5506 219020
rect 128357 219011 128415 219017
rect 128357 219008 128369 219011
rect 5500 218980 128369 219008
rect 5500 218968 5506 218980
rect 128357 218977 128369 218980
rect 128403 218977 128415 219011
rect 128357 218971 128415 218977
rect 4614 218900 4620 218952
rect 4672 218940 4678 218952
rect 128449 218943 128507 218949
rect 128449 218940 128461 218943
rect 4672 218912 128461 218940
rect 4672 218900 4678 218912
rect 128449 218909 128461 218912
rect 128495 218909 128507 218943
rect 224926 218940 224954 219320
rect 232958 219308 232964 219320
rect 233016 219308 233022 219360
rect 248322 219348 248328 219360
rect 248283 219320 248328 219348
rect 248322 219308 248328 219320
rect 248380 219308 248386 219360
rect 249426 219308 249432 219360
rect 249484 219348 249490 219360
rect 249484 219320 253934 219348
rect 249484 219308 249490 219320
rect 253906 219008 253934 219320
rect 260742 219308 260748 219360
rect 260800 219348 260806 219360
rect 260800 219320 267734 219348
rect 260800 219308 260806 219320
rect 267706 219076 267734 219320
rect 310974 219076 310980 219088
rect 267706 219048 310980 219076
rect 310974 219036 310980 219048
rect 311032 219036 311038 219088
rect 311526 219008 311532 219020
rect 253906 218980 311532 219008
rect 311526 218968 311532 218980
rect 311584 218968 311590 219020
rect 311802 218940 311808 218952
rect 224926 218912 311808 218940
rect 128449 218903 128507 218909
rect 311802 218900 311808 218912
rect 311860 218900 311866 218952
rect 8570 218832 8576 218884
rect 8628 218872 8634 218884
rect 78125 218875 78183 218881
rect 78125 218872 78137 218875
rect 8628 218844 78137 218872
rect 8628 218832 8634 218844
rect 78125 218841 78137 218844
rect 78171 218841 78183 218875
rect 78125 218835 78183 218841
rect 96065 218875 96123 218881
rect 96065 218841 96077 218875
rect 96111 218872 96123 218875
rect 310790 218872 310796 218884
rect 96111 218844 310796 218872
rect 96111 218841 96123 218844
rect 96065 218835 96123 218841
rect 310790 218832 310796 218844
rect 310848 218832 310854 218884
rect 8754 218764 8760 218816
rect 8812 218804 8818 218816
rect 22925 218807 22983 218813
rect 22925 218804 22937 218807
rect 8812 218776 22937 218804
rect 8812 218764 8818 218776
rect 22925 218773 22937 218776
rect 22971 218773 22983 218807
rect 22925 218767 22983 218773
rect 53745 218807 53803 218813
rect 53745 218773 53757 218807
rect 53791 218804 53803 218807
rect 483842 218804 483848 218816
rect 53791 218776 483848 218804
rect 53791 218773 53803 218776
rect 53745 218767 53803 218773
rect 483842 218764 483848 218776
rect 483900 218764 483906 218816
rect 9490 218696 9496 218748
rect 9548 218736 9554 218748
rect 232961 218739 233019 218745
rect 232961 218736 232973 218739
rect 9548 218708 232973 218736
rect 9548 218696 9554 218708
rect 232961 218705 232973 218708
rect 233007 218705 233019 218739
rect 232961 218699 233019 218705
rect 248325 218739 248383 218745
rect 248325 218705 248337 218739
rect 248371 218736 248383 218739
rect 310882 218736 310888 218748
rect 248371 218708 310888 218736
rect 248371 218705 248383 218708
rect 248325 218699 248383 218705
rect 310882 218696 310888 218708
rect 310940 218696 310946 218748
rect 6914 218628 6920 218680
rect 6972 218668 6978 218680
rect 17221 218671 17279 218677
rect 17221 218668 17233 218671
rect 6972 218640 17233 218668
rect 6972 218628 6978 218640
rect 17221 218637 17233 218640
rect 17267 218637 17279 218671
rect 17221 218631 17279 218637
rect 6730 218560 6736 218612
rect 6788 218600 6794 218612
rect 16209 218603 16267 218609
rect 16209 218600 16221 218603
rect 6788 218572 16221 218600
rect 6788 218560 6794 218572
rect 16209 218569 16221 218572
rect 16255 218569 16267 218603
rect 16209 218563 16267 218569
rect 5718 218492 5724 218544
rect 5776 218532 5782 218544
rect 12805 218535 12863 218541
rect 12805 218532 12817 218535
rect 5776 218504 12817 218532
rect 5776 218492 5782 218504
rect 12805 218501 12817 218504
rect 12851 218501 12863 218535
rect 12805 218495 12863 218501
rect 7282 218424 7288 218476
rect 7340 218464 7346 218476
rect 11793 218467 11851 218473
rect 11793 218464 11805 218467
rect 7340 218436 11805 218464
rect 7340 218424 7346 218436
rect 11793 218433 11805 218436
rect 11839 218433 11851 218467
rect 11793 218427 11851 218433
rect 114373 218263 114431 218269
rect 114373 218229 114385 218263
rect 114419 218260 114431 218263
rect 345845 218263 345903 218269
rect 345845 218260 345857 218263
rect 114419 218232 345857 218260
rect 114419 218229 114431 218232
rect 114373 218223 114431 218229
rect 345845 218229 345857 218232
rect 345891 218229 345903 218263
rect 345845 218223 345903 218229
rect 399478 218016 399484 218068
rect 399536 218056 399542 218068
rect 495434 218056 495440 218068
rect 399536 218028 495440 218056
rect 399536 218016 399542 218028
rect 495434 218016 495440 218028
rect 495492 218016 495498 218068
rect 9490 217716 9496 217728
rect 9451 217688 9496 217716
rect 9490 217676 9496 217688
rect 9548 217676 9554 217728
rect 3602 217608 3608 217660
rect 3660 217648 3666 217660
rect 310514 217648 310520 217660
rect 3660 217620 310520 217648
rect 3660 217608 3666 217620
rect 310514 217608 310520 217620
rect 310572 217608 310578 217660
rect 8386 217540 8392 217592
rect 8444 217580 8450 217592
rect 485406 217580 485412 217592
rect 8444 217552 485412 217580
rect 8444 217540 8450 217552
rect 485406 217540 485412 217552
rect 485464 217540 485470 217592
rect 7466 217472 7472 217524
rect 7524 217512 7530 217524
rect 496354 217512 496360 217524
rect 7524 217484 496360 217512
rect 7524 217472 7530 217484
rect 496354 217472 496360 217484
rect 496412 217472 496418 217524
rect 370961 216971 371019 216977
rect 370961 216968 370973 216971
rect 354646 216940 360194 216968
rect 312538 216792 312544 216844
rect 312596 216832 312602 216844
rect 354646 216832 354674 216940
rect 312596 216804 354674 216832
rect 360166 216832 360194 216940
rect 367066 216940 370973 216968
rect 367066 216832 367094 216940
rect 370961 216937 370973 216940
rect 371007 216937 371019 216971
rect 370961 216931 371019 216937
rect 371142 216928 371148 216980
rect 371200 216968 371206 216980
rect 371200 216940 379514 216968
rect 371200 216928 371206 216940
rect 370869 216903 370927 216909
rect 370869 216869 370881 216903
rect 370915 216900 370927 216903
rect 379486 216900 379514 216940
rect 428918 216900 428924 216912
rect 370915 216872 371556 216900
rect 379486 216872 428924 216900
rect 370915 216869 370927 216872
rect 370869 216863 370927 216869
rect 360166 216804 367094 216832
rect 370961 216835 371019 216841
rect 312596 216792 312602 216804
rect 370961 216801 370973 216835
rect 371007 216832 371019 216835
rect 371237 216835 371295 216841
rect 371237 216832 371249 216835
rect 371007 216804 371249 216832
rect 371007 216801 371019 216804
rect 370961 216795 371019 216801
rect 371237 216801 371249 216804
rect 371283 216801 371295 216835
rect 371237 216795 371295 216801
rect 313182 216724 313188 216776
rect 313240 216764 313246 216776
rect 370869 216767 370927 216773
rect 370869 216764 370881 216767
rect 313240 216736 370881 216764
rect 313240 216724 313246 216736
rect 370869 216733 370881 216736
rect 370915 216733 370927 216767
rect 371142 216764 371148 216776
rect 371103 216736 371148 216764
rect 370869 216727 370927 216733
rect 371142 216724 371148 216736
rect 371200 216724 371206 216776
rect 371418 216764 371424 216776
rect 371379 216736 371424 216764
rect 371418 216724 371424 216736
rect 371476 216724 371482 216776
rect 371528 216773 371556 216872
rect 428918 216860 428924 216872
rect 428976 216860 428982 216912
rect 371513 216767 371571 216773
rect 371513 216733 371525 216767
rect 371559 216733 371571 216767
rect 371513 216727 371571 216733
rect 340414 216656 340420 216708
rect 340472 216696 340478 216708
rect 371697 216699 371755 216705
rect 371697 216696 371709 216699
rect 340472 216668 371709 216696
rect 340472 216656 340478 216668
rect 371697 216665 371709 216668
rect 371743 216665 371755 216699
rect 371697 216659 371755 216665
rect 310057 210443 310115 210449
rect 310057 210409 310069 210443
rect 310103 210440 310115 210443
rect 310514 210440 310520 210452
rect 310103 210412 310520 210440
rect 310103 210409 310115 210412
rect 310057 210403 310115 210409
rect 310514 210400 310520 210412
rect 310572 210400 310578 210452
rect 3237 209559 3295 209565
rect 3237 209525 3249 209559
rect 3283 209556 3295 209559
rect 5994 209556 6000 209568
rect 3283 209528 6000 209556
rect 3283 209525 3295 209528
rect 3237 209519 3295 209525
rect 5994 209516 6000 209528
rect 6052 209516 6058 209568
rect 2866 205980 2872 206032
rect 2924 206020 2930 206032
rect 5626 206020 5632 206032
rect 2924 205992 5632 206020
rect 2924 205980 2930 205992
rect 5626 205980 5632 205992
rect 5684 205980 5690 206032
rect 8662 203872 8668 203924
rect 8720 203912 8726 203924
rect 9490 203912 9496 203924
rect 8720 203884 9496 203912
rect 8720 203872 8726 203884
rect 9490 203872 9496 203884
rect 9548 203872 9554 203924
rect 5626 203668 5632 203720
rect 5684 203708 5690 203720
rect 9309 203711 9367 203717
rect 9309 203708 9321 203711
rect 5684 203680 9321 203708
rect 5684 203668 5690 203680
rect 9309 203677 9321 203680
rect 9355 203677 9367 203711
rect 9309 203671 9367 203677
rect 331214 202784 331220 202836
rect 331272 202824 331278 202836
rect 467374 202824 467380 202836
rect 331272 202796 467380 202824
rect 331272 202784 331278 202796
rect 467374 202784 467380 202796
rect 467432 202784 467438 202836
rect 310057 202147 310115 202153
rect 310057 202113 310069 202147
rect 310103 202144 310115 202147
rect 311066 202144 311072 202156
rect 310103 202116 311072 202144
rect 310103 202113 310115 202116
rect 310057 202107 310115 202113
rect 311066 202104 311072 202116
rect 311124 202104 311130 202156
rect 311802 202008 311808 202020
rect 310348 201980 311808 202008
rect 310348 201949 310376 201980
rect 311802 201968 311808 201980
rect 311860 201968 311866 202020
rect 310333 201943 310391 201949
rect 310333 201909 310345 201943
rect 310379 201909 310391 201943
rect 310333 201903 310391 201909
rect 310517 201943 310575 201949
rect 310517 201909 310529 201943
rect 310563 201940 310575 201943
rect 331214 201940 331220 201952
rect 310563 201912 331220 201940
rect 310563 201909 310575 201912
rect 310517 201903 310575 201909
rect 331214 201900 331220 201912
rect 331272 201900 331278 201952
rect 313826 201424 313832 201476
rect 313884 201464 313890 201476
rect 495434 201464 495440 201476
rect 313884 201436 495440 201464
rect 313884 201424 313890 201436
rect 495434 201424 495440 201436
rect 495492 201424 495498 201476
rect 322198 200812 322204 200864
rect 322256 200852 322262 200864
rect 413741 200855 413799 200861
rect 413741 200852 413753 200855
rect 322256 200824 413753 200852
rect 322256 200812 322262 200824
rect 413741 200821 413753 200824
rect 413787 200821 413799 200855
rect 413741 200815 413799 200821
rect 483842 199968 483848 199980
rect 483803 199940 483848 199968
rect 483842 199928 483848 199940
rect 483900 199928 483906 199980
rect 3234 197752 3240 197804
rect 3292 197792 3298 197804
rect 7558 197792 7564 197804
rect 3292 197764 7564 197792
rect 3292 197752 3298 197764
rect 7558 197752 7564 197764
rect 7616 197752 7622 197804
rect 405918 197276 405924 197328
rect 405976 197316 405982 197328
rect 495434 197316 495440 197328
rect 405976 197288 495440 197316
rect 405976 197276 405982 197288
rect 495434 197276 495440 197288
rect 495492 197276 495498 197328
rect 349798 195372 349804 195424
rect 349856 195412 349862 195424
rect 450541 195415 450599 195421
rect 450541 195412 450553 195415
rect 349856 195384 450553 195412
rect 349856 195372 349862 195384
rect 450541 195381 450553 195384
rect 450587 195381 450599 195415
rect 450541 195375 450599 195381
rect 315758 194964 315764 195016
rect 315816 195004 315822 195016
rect 397457 195007 397515 195013
rect 397457 195004 397469 195007
rect 315816 194976 397469 195004
rect 315816 194964 315822 194976
rect 397457 194973 397469 194976
rect 397503 194973 397515 195007
rect 397457 194967 397515 194973
rect 472618 191836 472624 191888
rect 472676 191876 472682 191888
rect 495434 191876 495440 191888
rect 472676 191848 495440 191876
rect 472676 191836 472682 191848
rect 495434 191836 495440 191848
rect 495492 191836 495498 191888
rect 349798 187688 349804 187740
rect 349856 187728 349862 187740
rect 495434 187728 495440 187740
rect 349856 187700 495440 187728
rect 349856 187688 349862 187700
rect 495434 187688 495440 187700
rect 495492 187688 495498 187740
rect 310330 183948 310336 184000
rect 310388 183988 310394 184000
rect 310388 183960 316034 183988
rect 310388 183948 310394 183960
rect 311618 183784 311624 183796
rect 310440 183756 311624 183784
rect 310330 183648 310336 183660
rect 310291 183620 310336 183648
rect 310330 183608 310336 183620
rect 310388 183608 310394 183660
rect 310440 183657 310468 183756
rect 311618 183744 311624 183756
rect 311676 183744 311682 183796
rect 310790 183716 310796 183728
rect 310532 183688 310796 183716
rect 310532 183657 310560 183688
rect 310790 183676 310796 183688
rect 310848 183676 310854 183728
rect 316006 183716 316034 183960
rect 469858 183716 469864 183728
rect 316006 183688 469864 183716
rect 469858 183676 469864 183688
rect 469916 183676 469922 183728
rect 310425 183651 310483 183657
rect 310425 183617 310437 183651
rect 310471 183617 310483 183651
rect 310425 183611 310483 183617
rect 310517 183651 310575 183657
rect 310517 183617 310529 183651
rect 310563 183617 310575 183651
rect 310517 183611 310575 183617
rect 310698 183608 310704 183660
rect 310756 183648 310762 183660
rect 311802 183648 311808 183660
rect 310756 183620 311808 183648
rect 310756 183608 310762 183620
rect 311802 183608 311808 183620
rect 311860 183648 311866 183660
rect 311860 183620 316034 183648
rect 311860 183608 311866 183620
rect 310057 183583 310115 183589
rect 310057 183549 310069 183583
rect 310103 183580 310115 183583
rect 310606 183580 310612 183592
rect 310103 183552 310612 183580
rect 310103 183549 310115 183552
rect 310057 183543 310115 183549
rect 310606 183540 310612 183552
rect 310664 183540 310670 183592
rect 316006 183580 316034 183620
rect 453022 183580 453028 183592
rect 316006 183552 453028 183580
rect 453022 183540 453028 183552
rect 453080 183540 453086 183592
rect 3050 183404 3056 183456
rect 3108 183444 3114 183456
rect 6086 183444 6092 183456
rect 3108 183416 6092 183444
rect 3108 183404 3114 183416
rect 6086 183404 6092 183416
rect 6144 183404 6150 183456
rect 406378 179772 406384 179784
rect 406339 179744 406384 179772
rect 406378 179732 406384 179744
rect 406436 179732 406442 179784
rect 407577 179775 407635 179781
rect 407577 179772 407589 179775
rect 406856 179744 407589 179772
rect 406856 179645 406884 179744
rect 407577 179741 407589 179744
rect 407623 179741 407635 179775
rect 407577 179735 407635 179741
rect 406841 179639 406899 179645
rect 406841 179605 406853 179639
rect 406887 179605 406899 179639
rect 407390 179636 407396 179648
rect 407351 179608 407396 179636
rect 406841 179599 406899 179605
rect 407390 179596 407396 179608
rect 407448 179596 407454 179648
rect 3326 178848 3332 178900
rect 3384 178888 3390 178900
rect 3970 178888 3976 178900
rect 3384 178860 3976 178888
rect 3384 178848 3390 178860
rect 3970 178848 3976 178860
rect 4028 178848 4034 178900
rect 310698 178508 310704 178560
rect 310756 178548 310762 178560
rect 346854 178548 346860 178560
rect 310756 178520 346860 178548
rect 310756 178508 310762 178520
rect 346854 178508 346860 178520
rect 346912 178508 346918 178560
rect 310149 178347 310207 178353
rect 310149 178313 310161 178347
rect 310195 178344 310207 178347
rect 310882 178344 310888 178356
rect 310195 178316 310888 178344
rect 310195 178313 310207 178316
rect 310149 178307 310207 178313
rect 310882 178304 310888 178316
rect 310940 178304 310946 178356
rect 310514 178276 310520 178288
rect 310348 178248 310520 178276
rect 310348 178217 310376 178248
rect 310514 178236 310520 178248
rect 310572 178276 310578 178288
rect 311526 178276 311532 178288
rect 310572 178248 311532 178276
rect 310572 178236 310578 178248
rect 311526 178236 311532 178248
rect 311584 178236 311590 178288
rect 311866 178248 316034 178276
rect 310333 178211 310391 178217
rect 310333 178177 310345 178211
rect 310379 178177 310391 178211
rect 310333 178171 310391 178177
rect 310422 178168 310428 178220
rect 310480 178208 310486 178220
rect 311866 178208 311894 178248
rect 310480 178180 311894 178208
rect 316006 178208 316034 178248
rect 407390 178208 407396 178220
rect 316006 178180 407396 178208
rect 310480 178168 310486 178180
rect 407390 178168 407396 178180
rect 407448 178168 407454 178220
rect 310698 178140 310704 178152
rect 310659 178112 310704 178140
rect 310698 178100 310704 178112
rect 310756 178100 310762 178152
rect 310609 178075 310667 178081
rect 310609 178041 310621 178075
rect 310655 178072 310667 178075
rect 310790 178072 310796 178084
rect 310655 178044 310796 178072
rect 310655 178041 310667 178044
rect 310609 178035 310667 178041
rect 310790 178032 310796 178044
rect 310848 178032 310854 178084
rect 310238 176168 310244 176180
rect 310199 176140 310244 176168
rect 310238 176128 310244 176140
rect 310296 176128 310302 176180
rect 336182 176168 336188 176180
rect 336143 176140 336188 176168
rect 336182 176128 336188 176140
rect 336240 176128 336246 176180
rect 336550 176168 336556 176180
rect 336511 176140 336556 176168
rect 336550 176128 336556 176140
rect 336608 176128 336614 176180
rect 336090 176100 336096 176112
rect 336051 176072 336096 176100
rect 336090 176060 336096 176072
rect 336148 176060 336154 176112
rect 310057 176035 310115 176041
rect 310057 176001 310069 176035
rect 310103 176032 310115 176035
rect 310698 176032 310704 176044
rect 310103 176004 310704 176032
rect 310103 176001 310115 176004
rect 310057 175995 310115 176001
rect 310698 175992 310704 176004
rect 310756 176032 310762 176044
rect 310974 176032 310980 176044
rect 310756 176004 310980 176032
rect 310756 175992 310762 176004
rect 310974 175992 310980 176004
rect 311032 175992 311038 176044
rect 335906 175964 335912 175976
rect 335867 175936 335912 175964
rect 335906 175924 335912 175936
rect 335964 175964 335970 175976
rect 337013 175967 337071 175973
rect 337013 175964 337025 175967
rect 335964 175936 337025 175964
rect 335964 175924 335970 175936
rect 337013 175933 337025 175936
rect 337059 175933 337071 175967
rect 337013 175927 337071 175933
rect 337470 175828 337476 175840
rect 337431 175800 337476 175828
rect 337470 175788 337476 175800
rect 337528 175788 337534 175840
rect 310238 175584 310244 175636
rect 310296 175624 310302 175636
rect 419534 175624 419540 175636
rect 310296 175596 419540 175624
rect 310296 175584 310302 175596
rect 419534 175584 419540 175596
rect 419592 175584 419598 175636
rect 324958 175176 324964 175228
rect 325016 175216 325022 175228
rect 495434 175216 495440 175228
rect 325016 175188 495440 175216
rect 325016 175176 325022 175188
rect 495434 175176 495440 175188
rect 495492 175176 495498 175228
rect 3326 170144 3332 170196
rect 3384 170184 3390 170196
rect 3605 170187 3663 170193
rect 3605 170184 3617 170187
rect 3384 170156 3617 170184
rect 3384 170144 3390 170156
rect 3605 170153 3617 170156
rect 3651 170153 3663 170187
rect 3605 170147 3663 170153
rect 4985 170051 5043 170057
rect 4985 170017 4997 170051
rect 5031 170048 5043 170051
rect 5166 170048 5172 170060
rect 5031 170020 5172 170048
rect 5031 170017 5043 170020
rect 4985 170011 5043 170017
rect 5166 170008 5172 170020
rect 5224 170008 5230 170060
rect 4729 169983 4787 169989
rect 4729 169949 4741 169983
rect 4775 169980 4787 169983
rect 5074 169980 5080 169992
rect 4775 169952 5080 169980
rect 4775 169949 4787 169952
rect 4729 169943 4787 169949
rect 5074 169940 5080 169952
rect 5132 169940 5138 169992
rect 3970 169804 3976 169856
rect 4028 169844 4034 169856
rect 7374 169844 7380 169856
rect 4028 169816 7380 169844
rect 4028 169804 4034 169816
rect 7374 169804 7380 169816
rect 7432 169804 7438 169856
rect 380618 161984 380624 162036
rect 380676 162024 380682 162036
rect 380713 162027 380771 162033
rect 380713 162024 380725 162027
rect 380676 161996 380725 162024
rect 380676 161984 380682 161996
rect 380713 161993 380725 161996
rect 380759 161993 380771 162027
rect 381078 162024 381084 162036
rect 381039 161996 381084 162024
rect 380713 161987 380771 161993
rect 381078 161984 381084 161996
rect 381136 161984 381142 162036
rect 424042 162024 424048 162036
rect 385604 161996 424048 162024
rect 378778 161916 378784 161968
rect 378836 161956 378842 161968
rect 385405 161959 385463 161965
rect 385405 161956 385417 161959
rect 378836 161928 385417 161956
rect 378836 161916 378842 161928
rect 385405 161925 385417 161928
rect 385451 161925 385463 161959
rect 385405 161919 385463 161925
rect 385604 161900 385632 161996
rect 424042 161984 424048 161996
rect 424100 161984 424106 162036
rect 470502 161956 470508 161968
rect 385788 161928 470508 161956
rect 385788 161900 385816 161928
rect 470502 161916 470508 161928
rect 470560 161916 470566 161968
rect 385034 161888 385040 161900
rect 384995 161860 385040 161888
rect 385034 161848 385040 161860
rect 385092 161848 385098 161900
rect 385218 161888 385224 161900
rect 385179 161860 385224 161888
rect 385218 161848 385224 161860
rect 385276 161848 385282 161900
rect 385586 161888 385592 161900
rect 385499 161860 385592 161888
rect 385586 161848 385592 161860
rect 385644 161848 385650 161900
rect 385770 161888 385776 161900
rect 385683 161860 385776 161888
rect 385770 161848 385776 161860
rect 385828 161848 385834 161900
rect 419074 161888 419080 161900
rect 393286 161860 419080 161888
rect 380158 161780 380164 161832
rect 380216 161820 380222 161832
rect 381173 161823 381231 161829
rect 381173 161820 381185 161823
rect 380216 161792 381185 161820
rect 380216 161780 380222 161792
rect 381173 161789 381185 161792
rect 381219 161789 381231 161823
rect 381173 161783 381231 161789
rect 381357 161823 381415 161829
rect 381357 161789 381369 161823
rect 381403 161820 381415 161823
rect 382182 161820 382188 161832
rect 381403 161792 382188 161820
rect 381403 161789 381415 161792
rect 381357 161783 381415 161789
rect 382182 161780 382188 161792
rect 382240 161820 382246 161832
rect 382240 161792 383654 161820
rect 382240 161780 382246 161792
rect 383626 161752 383654 161792
rect 393286 161752 393314 161860
rect 419074 161848 419080 161860
rect 419132 161848 419138 161900
rect 383626 161724 393314 161752
rect 414842 161684 414848 161696
rect 414803 161656 414848 161684
rect 414842 161644 414848 161656
rect 414900 161644 414906 161696
rect 465997 161687 466055 161693
rect 465997 161684 466009 161687
rect 451246 161656 466009 161684
rect 315942 161440 315948 161492
rect 316000 161480 316006 161492
rect 451246 161480 451274 161656
rect 465997 161653 466009 161656
rect 466043 161653 466055 161687
rect 465997 161647 466055 161653
rect 316000 161452 451274 161480
rect 316000 161440 316006 161452
rect 3326 161100 3332 161152
rect 3384 161140 3390 161152
rect 6454 161140 6460 161152
rect 3384 161112 6460 161140
rect 3384 161100 3390 161112
rect 6454 161100 6460 161112
rect 6512 161100 6518 161152
rect 8113 157131 8171 157137
rect 8113 157097 8125 157131
rect 8159 157128 8171 157131
rect 9122 157128 9128 157140
rect 8159 157100 9128 157128
rect 8159 157097 8171 157100
rect 8113 157091 8171 157097
rect 9122 157088 9128 157100
rect 9180 157088 9186 157140
rect 484210 157128 484216 157140
rect 484171 157100 484216 157128
rect 484210 157088 484216 157100
rect 484268 157088 484274 157140
rect 3142 157020 3148 157072
rect 3200 157060 3206 157072
rect 6362 157060 6368 157072
rect 3200 157032 6368 157060
rect 3200 157020 3206 157032
rect 6362 157020 6368 157032
rect 6420 157020 6426 157072
rect 8205 156927 8263 156933
rect 8205 156893 8217 156927
rect 8251 156924 8263 156927
rect 8938 156924 8944 156936
rect 8251 156896 8944 156924
rect 8251 156893 8263 156896
rect 8205 156887 8263 156893
rect 8938 156884 8944 156896
rect 8996 156884 9002 156936
rect 321462 152640 321468 152652
rect 321423 152612 321468 152640
rect 321462 152600 321468 152612
rect 321520 152600 321526 152652
rect 323578 152640 323584 152652
rect 323539 152612 323584 152640
rect 323578 152600 323584 152612
rect 323636 152640 323642 152652
rect 323636 152612 325694 152640
rect 323636 152600 323642 152612
rect 325666 152572 325694 152612
rect 429194 152572 429200 152584
rect 325666 152544 429200 152572
rect 429194 152532 429200 152544
rect 429252 152532 429258 152584
rect 322017 152439 322075 152445
rect 322017 152405 322029 152439
rect 322063 152436 322075 152439
rect 322477 152439 322535 152445
rect 322063 152408 322428 152436
rect 322063 152405 322075 152408
rect 322017 152399 322075 152405
rect 322293 152167 322351 152173
rect 322293 152164 322305 152167
rect 321756 152136 322305 152164
rect 321756 152105 321784 152136
rect 322293 152133 322305 152136
rect 322339 152133 322351 152167
rect 322293 152127 322351 152133
rect 321649 152099 321707 152105
rect 321649 152065 321661 152099
rect 321695 152065 321707 152099
rect 321649 152059 321707 152065
rect 321741 152099 321799 152105
rect 321741 152065 321753 152099
rect 321787 152065 321799 152099
rect 321741 152059 321799 152065
rect 322017 152099 322075 152105
rect 322017 152065 322029 152099
rect 322063 152096 322075 152099
rect 322400 152096 322428 152408
rect 322477 152405 322489 152439
rect 322523 152436 322535 152439
rect 323029 152439 323087 152445
rect 323029 152436 323041 152439
rect 322523 152408 323041 152436
rect 322523 152405 322535 152408
rect 322477 152399 322535 152405
rect 323029 152405 323041 152408
rect 323075 152405 323087 152439
rect 323029 152399 323087 152405
rect 322063 152068 322428 152096
rect 322063 152065 322075 152068
rect 322017 152059 322075 152065
rect 321664 151972 321692 152059
rect 425698 152056 425704 152108
rect 425756 152096 425762 152108
rect 427265 152099 427323 152105
rect 427265 152096 427277 152099
rect 425756 152068 427277 152096
rect 425756 152056 425762 152068
rect 427265 152065 427277 152068
rect 427311 152065 427323 152099
rect 427265 152059 427323 152065
rect 321922 152028 321928 152040
rect 321883 152000 321928 152028
rect 321922 151988 321928 152000
rect 321980 151988 321986 152040
rect 417510 152028 417516 152040
rect 325666 152000 417516 152028
rect 321646 151960 321652 151972
rect 321559 151932 321652 151960
rect 321646 151920 321652 151932
rect 321704 151960 321710 151972
rect 325666 151960 325694 152000
rect 417510 151988 417516 152000
rect 417568 151988 417574 152040
rect 321704 151932 325694 151960
rect 321704 151920 321710 151932
rect 321370 151852 321376 151904
rect 321428 151892 321434 151904
rect 321465 151895 321523 151901
rect 321465 151892 321477 151895
rect 321428 151864 321477 151892
rect 321428 151852 321434 151864
rect 321465 151861 321477 151864
rect 321511 151861 321523 151895
rect 321465 151855 321523 151861
rect 357342 148220 357348 148232
rect 357303 148192 357348 148220
rect 357342 148180 357348 148192
rect 357400 148180 357406 148232
rect 315206 147500 315212 147552
rect 315264 147540 315270 147552
rect 315485 147543 315543 147549
rect 315485 147540 315497 147543
rect 315264 147512 315497 147540
rect 315264 147500 315270 147512
rect 315485 147509 315497 147512
rect 315531 147509 315543 147543
rect 315485 147503 315543 147509
rect 486970 146888 486976 146940
rect 487028 146928 487034 146940
rect 495526 146928 495532 146940
rect 487028 146900 495532 146928
rect 487028 146888 487034 146900
rect 495526 146888 495532 146900
rect 495584 146888 495590 146940
rect 9493 145367 9551 145373
rect 9493 145333 9505 145367
rect 9539 145364 9551 145367
rect 9539 145336 9628 145364
rect 9539 145333 9551 145336
rect 9493 145327 9551 145333
rect 9600 145169 9628 145336
rect 9585 145163 9643 145169
rect 9585 145129 9597 145163
rect 9631 145129 9643 145163
rect 9585 145123 9643 145129
rect 418154 143488 418160 143540
rect 418212 143528 418218 143540
rect 418798 143528 418804 143540
rect 418212 143500 418804 143528
rect 418212 143488 418218 143500
rect 418798 143488 418804 143500
rect 418856 143528 418862 143540
rect 495434 143528 495440 143540
rect 418856 143500 495440 143528
rect 418856 143488 418862 143500
rect 495434 143488 495440 143500
rect 495492 143488 495498 143540
rect 389358 143188 389364 143200
rect 389319 143160 389364 143188
rect 389358 143148 389364 143160
rect 389416 143148 389422 143200
rect 316586 142808 316592 142860
rect 316644 142848 316650 142860
rect 418154 142848 418160 142860
rect 316644 142820 418160 142848
rect 316644 142808 316650 142820
rect 418154 142808 418160 142820
rect 418212 142808 418218 142860
rect 361482 142740 361488 142792
rect 361540 142780 361546 142792
rect 454957 142783 455015 142789
rect 454957 142780 454969 142783
rect 361540 142752 454969 142780
rect 361540 142740 361546 142752
rect 454957 142749 454969 142752
rect 455003 142749 455015 142783
rect 454957 142743 455015 142749
rect 9766 142304 9772 142316
rect 9727 142276 9772 142304
rect 9766 142264 9772 142276
rect 9824 142264 9830 142316
rect 9585 142171 9643 142177
rect 9585 142137 9597 142171
rect 9631 142168 9643 142171
rect 9766 142168 9772 142180
rect 9631 142140 9772 142168
rect 9631 142137 9643 142140
rect 9585 142131 9643 142137
rect 9766 142128 9772 142140
rect 9824 142128 9830 142180
rect 313826 142128 313832 142180
rect 313884 142168 313890 142180
rect 457717 142171 457775 142177
rect 457717 142168 457729 142171
rect 313884 142140 457729 142168
rect 313884 142128 313890 142140
rect 457717 142137 457729 142140
rect 457763 142137 457775 142171
rect 457717 142131 457775 142137
rect 416130 140604 416136 140616
rect 416043 140576 416136 140604
rect 416130 140564 416136 140576
rect 416188 140604 416194 140616
rect 451642 140604 451648 140616
rect 416188 140576 451648 140604
rect 416188 140564 416194 140576
rect 451642 140564 451648 140576
rect 451700 140564 451706 140616
rect 416406 140545 416412 140548
rect 416400 140499 416412 140545
rect 416464 140536 416470 140548
rect 416464 140508 416500 140536
rect 416406 140496 416412 140499
rect 416464 140496 416470 140508
rect 417418 140428 417424 140480
rect 417476 140468 417482 140480
rect 417513 140471 417571 140477
rect 417513 140468 417525 140471
rect 417476 140440 417525 140468
rect 417476 140428 417482 140440
rect 417513 140437 417525 140440
rect 417559 140468 417571 140471
rect 473630 140468 473636 140480
rect 417559 140440 473636 140468
rect 417559 140437 417571 140440
rect 417513 140431 417571 140437
rect 473630 140428 473636 140440
rect 473688 140428 473694 140480
rect 3326 138932 3332 138984
rect 3384 138972 3390 138984
rect 6546 138972 6552 138984
rect 3384 138944 6552 138972
rect 3384 138932 3390 138944
rect 6546 138932 6552 138944
rect 6604 138932 6610 138984
rect 8386 136416 8392 136468
rect 8444 136456 8450 136468
rect 9122 136456 9128 136468
rect 8444 136428 9128 136456
rect 8444 136416 8450 136428
rect 9122 136416 9128 136428
rect 9180 136456 9186 136468
rect 9401 136459 9459 136465
rect 9401 136456 9413 136459
rect 9180 136428 9413 136456
rect 9180 136416 9186 136428
rect 9401 136425 9413 136428
rect 9447 136425 9459 136459
rect 9401 136419 9459 136425
rect 7469 136391 7527 136397
rect 7469 136357 7481 136391
rect 7515 136388 7527 136391
rect 9769 136391 9827 136397
rect 9769 136388 9781 136391
rect 7515 136360 9781 136388
rect 7515 136357 7527 136360
rect 7469 136351 7527 136357
rect 9769 136357 9781 136360
rect 9815 136357 9827 136391
rect 9769 136351 9827 136357
rect 8478 136212 8484 136264
rect 8536 136252 8542 136264
rect 8938 136252 8944 136264
rect 8536 136224 8944 136252
rect 8536 136212 8542 136224
rect 8938 136212 8944 136224
rect 8996 136252 9002 136264
rect 9309 136255 9367 136261
rect 9309 136252 9321 136255
rect 8996 136224 9321 136252
rect 8996 136212 9002 136224
rect 9309 136221 9321 136224
rect 9355 136221 9367 136255
rect 9309 136215 9367 136221
rect 7285 135371 7343 135377
rect 7285 135337 7297 135371
rect 7331 135368 7343 135371
rect 7469 135371 7527 135377
rect 7469 135368 7481 135371
rect 7331 135340 7481 135368
rect 7331 135337 7343 135340
rect 7285 135331 7343 135337
rect 7469 135337 7481 135340
rect 7515 135337 7527 135371
rect 7469 135331 7527 135337
rect 8570 133084 8576 133136
rect 8628 133124 8634 133136
rect 8757 133127 8815 133133
rect 8757 133124 8769 133127
rect 8628 133096 8769 133124
rect 8628 133084 8634 133096
rect 8757 133093 8769 133096
rect 8803 133093 8815 133127
rect 8757 133087 8815 133093
rect 9030 133056 9036 133068
rect 8956 133028 9036 133056
rect 8956 132997 8984 133028
rect 9030 133016 9036 133028
rect 9088 133016 9094 133068
rect 9214 133056 9220 133068
rect 9175 133028 9220 133056
rect 9214 133016 9220 133028
rect 9272 133016 9278 133068
rect 9398 133056 9404 133068
rect 9324 133028 9404 133056
rect 9324 132997 9352 133028
rect 9398 133016 9404 133028
rect 9456 133016 9462 133068
rect 8941 132991 8999 132997
rect 8941 132957 8953 132991
rect 8987 132957 8999 132991
rect 8941 132951 8999 132957
rect 9125 132991 9183 132997
rect 9125 132957 9137 132991
rect 9171 132957 9183 132991
rect 9125 132951 9183 132957
rect 9310 132991 9368 132997
rect 9310 132957 9322 132991
rect 9356 132957 9368 132991
rect 9490 132988 9496 133000
rect 9451 132960 9496 132988
rect 9310 132951 9368 132957
rect 9140 132864 9168 132951
rect 9490 132948 9496 132960
rect 9548 132948 9554 133000
rect 355965 132991 356023 132997
rect 355965 132957 355977 132991
rect 356011 132988 356023 132991
rect 369302 132988 369308 133000
rect 356011 132960 369308 132988
rect 356011 132957 356023 132960
rect 355965 132951 356023 132957
rect 369302 132948 369308 132960
rect 369360 132948 369366 133000
rect 9398 132880 9404 132932
rect 9456 132920 9462 132932
rect 9858 132920 9864 132932
rect 9456 132892 9864 132920
rect 9456 132880 9462 132892
rect 9858 132880 9864 132892
rect 9916 132880 9922 132932
rect 9122 132812 9128 132864
rect 9180 132812 9186 132864
rect 319438 130364 319444 130416
rect 319496 130404 319502 130416
rect 482646 130404 482652 130416
rect 319496 130376 482652 130404
rect 319496 130364 319502 130376
rect 482646 130364 482652 130376
rect 482704 130364 482710 130416
rect 5350 129820 5356 129872
rect 5408 129860 5414 129872
rect 8202 129860 8208 129872
rect 5408 129832 8208 129860
rect 5408 129820 5414 129832
rect 8202 129820 8208 129832
rect 8260 129820 8266 129872
rect 356701 128639 356759 128645
rect 356701 128605 356713 128639
rect 356747 128636 356759 128639
rect 356790 128636 356796 128648
rect 356747 128608 356796 128636
rect 356747 128605 356759 128608
rect 356701 128599 356759 128605
rect 356790 128596 356796 128608
rect 356848 128596 356854 128648
rect 4522 127548 4528 127560
rect 4483 127520 4528 127548
rect 4522 127508 4528 127520
rect 4580 127508 4586 127560
rect 4709 127415 4767 127421
rect 4709 127381 4721 127415
rect 4755 127412 4767 127415
rect 5074 127412 5080 127424
rect 4755 127384 5080 127412
rect 4755 127381 4767 127384
rect 4709 127375 4767 127381
rect 5074 127372 5080 127384
rect 5132 127372 5138 127424
rect 363598 126420 363604 126472
rect 363656 126460 363662 126472
rect 383657 126463 383715 126469
rect 383657 126460 383669 126463
rect 363656 126432 383669 126460
rect 363656 126420 363662 126432
rect 383657 126429 383669 126432
rect 383703 126429 383715 126463
rect 383657 126423 383715 126429
rect 312262 126284 312268 126336
rect 312320 126324 312326 126336
rect 426618 126324 426624 126336
rect 312320 126296 426624 126324
rect 312320 126284 312326 126296
rect 426618 126284 426624 126296
rect 426676 126284 426682 126336
rect 477770 126120 477776 126132
rect 477731 126092 477776 126120
rect 477770 126080 477776 126092
rect 477828 126080 477834 126132
rect 311526 125944 311532 125996
rect 311584 125984 311590 125996
rect 312170 125984 312176 125996
rect 311584 125956 312176 125984
rect 311584 125944 311590 125956
rect 312170 125944 312176 125956
rect 312228 125944 312234 125996
rect 477678 125984 477684 125996
rect 477639 125956 477684 125984
rect 477678 125944 477684 125956
rect 477736 125944 477742 125996
rect 3970 125536 3976 125588
rect 4028 125576 4034 125588
rect 5350 125576 5356 125588
rect 4028 125548 5356 125576
rect 4028 125536 4034 125548
rect 5350 125536 5356 125548
rect 5408 125536 5414 125588
rect 428918 124896 428924 124908
rect 428879 124868 428924 124896
rect 428918 124856 428924 124868
rect 428976 124856 428982 124908
rect 429194 124896 429200 124908
rect 429155 124868 429200 124896
rect 429194 124856 429200 124868
rect 429252 124856 429258 124908
rect 429286 124856 429292 124908
rect 429344 124896 429350 124908
rect 429344 124868 429389 124896
rect 429344 124856 429350 124868
rect 384298 124720 384304 124772
rect 384356 124760 384362 124772
rect 429473 124763 429531 124769
rect 429473 124760 429485 124763
rect 384356 124732 429485 124760
rect 384356 124720 384362 124732
rect 429473 124729 429485 124732
rect 429519 124729 429531 124763
rect 429473 124723 429531 124729
rect 360838 124652 360844 124704
rect 360896 124692 360902 124704
rect 429013 124695 429071 124701
rect 429013 124692 429025 124695
rect 360896 124664 429025 124692
rect 360896 124652 360902 124664
rect 429013 124661 429025 124664
rect 429059 124661 429071 124695
rect 429013 124655 429071 124661
rect 310241 123607 310299 123613
rect 310241 123573 310253 123607
rect 310287 123604 310299 123607
rect 331858 123604 331864 123616
rect 310287 123576 331864 123604
rect 310287 123573 310299 123576
rect 310241 123567 310299 123573
rect 331858 123564 331864 123576
rect 331916 123564 331922 123616
rect 366818 123400 366824 123412
rect 366779 123372 366824 123400
rect 366818 123360 366824 123372
rect 366876 123360 366882 123412
rect 366726 123264 366732 123276
rect 366687 123236 366732 123264
rect 366726 123224 366732 123236
rect 366784 123224 366790 123276
rect 367002 123196 367008 123208
rect 366963 123168 367008 123196
rect 367002 123156 367008 123168
rect 367060 123156 367066 123208
rect 367094 123156 367100 123208
rect 367152 123196 367158 123208
rect 367152 123168 367197 123196
rect 367152 123156 367158 123168
rect 318150 123020 318156 123072
rect 318208 123060 318214 123072
rect 367281 123063 367339 123069
rect 367281 123060 367293 123063
rect 318208 123032 367293 123060
rect 318208 123020 318214 123032
rect 367281 123029 367293 123032
rect 367327 123029 367339 123063
rect 367281 123023 367339 123029
rect 9122 121864 9128 121916
rect 9180 121904 9186 121916
rect 385586 121904 385592 121916
rect 9180 121876 385592 121904
rect 9180 121864 9186 121876
rect 385586 121864 385592 121876
rect 385644 121864 385650 121916
rect 4062 121796 4068 121848
rect 4120 121836 4126 121848
rect 321646 121836 321652 121848
rect 4120 121808 321652 121836
rect 4120 121796 4126 121808
rect 321646 121796 321652 121808
rect 321704 121796 321710 121848
rect 9490 121728 9496 121780
rect 9548 121768 9554 121780
rect 311802 121768 311808 121780
rect 9548 121740 311808 121768
rect 9548 121728 9554 121740
rect 311802 121728 311808 121740
rect 311860 121728 311866 121780
rect 2774 121116 2780 121168
rect 2832 121156 2838 121168
rect 5258 121156 5264 121168
rect 2832 121128 5264 121156
rect 2832 121116 2838 121128
rect 5258 121116 5264 121128
rect 5316 121116 5322 121168
rect 299661 120887 299719 120893
rect 299661 120853 299673 120887
rect 299707 120884 299719 120887
rect 311986 120884 311992 120896
rect 299707 120856 311992 120884
rect 299707 120853 299719 120856
rect 299661 120847 299719 120853
rect 311986 120844 311992 120856
rect 312044 120844 312050 120896
rect 7190 120776 7196 120828
rect 7248 120816 7254 120828
rect 248877 120819 248935 120825
rect 7248 120788 20760 120816
rect 7248 120776 7254 120788
rect 20732 120760 20760 120788
rect 248877 120785 248889 120819
rect 248923 120816 248935 120819
rect 311066 120816 311072 120828
rect 248923 120788 311072 120816
rect 248923 120785 248935 120788
rect 248877 120779 248935 120785
rect 311066 120776 311072 120788
rect 311124 120776 311130 120828
rect 20714 120708 20720 120760
rect 20772 120708 20778 120760
rect 128998 120748 129004 120760
rect 26206 120720 129004 120748
rect 7098 120572 7104 120624
rect 7156 120612 7162 120624
rect 26206 120612 26234 120720
rect 128998 120708 129004 120720
rect 129056 120708 129062 120760
rect 216122 120708 216128 120760
rect 216180 120748 216186 120760
rect 310606 120748 310612 120760
rect 216180 120720 310612 120748
rect 216180 120708 216186 120720
rect 310606 120708 310612 120720
rect 310664 120708 310670 120760
rect 248874 120680 248880 120692
rect 248835 120652 248880 120680
rect 248874 120640 248880 120652
rect 248932 120640 248938 120692
rect 299658 120680 299664 120692
rect 299619 120652 299664 120680
rect 299658 120640 299664 120652
rect 299716 120640 299722 120692
rect 7156 120584 26234 120612
rect 7156 120572 7162 120584
rect 7006 120096 7012 120148
rect 7064 120136 7070 120148
rect 221826 120136 221832 120148
rect 7064 120108 221832 120136
rect 7064 120096 7070 120108
rect 221826 120096 221832 120108
rect 221884 120096 221890 120148
rect 239585 120071 239643 120077
rect 239585 120037 239597 120071
rect 239631 120068 239643 120071
rect 412082 120068 412088 120080
rect 239631 120040 412088 120068
rect 239631 120037 239643 120040
rect 239585 120031 239643 120037
rect 412082 120028 412088 120040
rect 412140 120028 412146 120080
rect 5718 119960 5724 120012
rect 5776 120000 5782 120012
rect 289817 120003 289875 120009
rect 289817 120000 289829 120003
rect 5776 119972 289829 120000
rect 5776 119960 5782 119972
rect 289817 119969 289829 119972
rect 289863 119969 289875 120003
rect 289817 119963 289875 119969
rect 289909 120003 289967 120009
rect 289909 119969 289921 120003
rect 289955 120000 289967 120003
rect 291841 120003 291899 120009
rect 291841 120000 291853 120003
rect 289955 119972 291853 120000
rect 289955 119969 289967 119972
rect 289909 119963 289967 119969
rect 291841 119969 291853 119972
rect 291887 119969 291899 120003
rect 291841 119963 291899 119969
rect 291933 120003 291991 120009
rect 291933 119969 291945 120003
rect 291979 120000 291991 120003
rect 477678 120000 477684 120012
rect 291979 119972 477684 120000
rect 291979 119969 291991 119972
rect 291933 119963 291991 119969
rect 477678 119960 477684 119972
rect 477736 119960 477742 120012
rect 156601 119935 156659 119941
rect 156601 119901 156613 119935
rect 156647 119932 156659 119935
rect 166261 119935 166319 119941
rect 166261 119932 166273 119935
rect 156647 119904 166273 119932
rect 156647 119901 156659 119904
rect 156601 119895 156659 119901
rect 166261 119901 166273 119904
rect 166307 119901 166319 119935
rect 166261 119895 166319 119901
rect 233881 119935 233939 119941
rect 233881 119901 233893 119935
rect 233927 119932 233939 119935
rect 239217 119935 239275 119941
rect 239217 119932 239229 119935
rect 233927 119904 239229 119932
rect 233927 119901 233939 119904
rect 233881 119895 233939 119901
rect 239217 119901 239229 119904
rect 239263 119901 239275 119935
rect 239217 119895 239275 119901
rect 239309 119935 239367 119941
rect 239309 119901 239321 119935
rect 239355 119932 239367 119935
rect 451550 119932 451556 119944
rect 239355 119904 451556 119932
rect 239355 119901 239367 119904
rect 239309 119895 239367 119901
rect 451550 119892 451556 119904
rect 451608 119892 451614 119944
rect 80977 119867 81035 119873
rect 80977 119833 80989 119867
rect 81023 119864 81035 119867
rect 311158 119864 311164 119876
rect 81023 119836 311164 119864
rect 81023 119833 81035 119836
rect 80977 119827 81035 119833
rect 311158 119824 311164 119836
rect 311216 119824 311222 119876
rect 75733 119799 75791 119805
rect 75733 119765 75745 119799
rect 75779 119796 75791 119799
rect 307665 119799 307723 119805
rect 307665 119796 307677 119799
rect 75779 119768 307677 119796
rect 75779 119765 75791 119768
rect 75733 119759 75791 119765
rect 307665 119765 307677 119768
rect 307711 119765 307723 119799
rect 307665 119759 307723 119765
rect 307772 119768 316034 119796
rect 258629 119731 258687 119737
rect 258629 119697 258641 119731
rect 258675 119728 258687 119731
rect 290001 119731 290059 119737
rect 290001 119728 290013 119731
rect 258675 119700 290013 119728
rect 258675 119697 258687 119700
rect 258629 119691 258687 119697
rect 290001 119697 290013 119700
rect 290047 119697 290059 119731
rect 290001 119691 290059 119697
rect 290737 119731 290795 119737
rect 290737 119697 290749 119731
rect 290783 119728 290795 119731
rect 307772 119728 307800 119768
rect 290783 119700 307800 119728
rect 308217 119731 308275 119737
rect 290783 119697 290795 119700
rect 290737 119691 290795 119697
rect 308217 119697 308229 119731
rect 308263 119728 308275 119731
rect 311342 119728 311348 119740
rect 308263 119700 311348 119728
rect 308263 119697 308275 119700
rect 308217 119691 308275 119697
rect 311342 119688 311348 119700
rect 311400 119688 311406 119740
rect 316006 119728 316034 119768
rect 342070 119728 342076 119740
rect 316006 119700 342076 119728
rect 342070 119688 342076 119700
rect 342128 119688 342134 119740
rect 216582 119620 216588 119672
rect 216640 119660 216646 119672
rect 233881 119663 233939 119669
rect 233881 119660 233893 119663
rect 216640 119632 233893 119660
rect 216640 119620 216646 119632
rect 233881 119629 233893 119632
rect 233927 119629 233939 119663
rect 233881 119623 233939 119629
rect 248509 119663 248567 119669
rect 248509 119629 248521 119663
rect 248555 119660 248567 119663
rect 253934 119660 253940 119672
rect 248555 119632 253940 119660
rect 248555 119629 248567 119632
rect 248509 119623 248567 119629
rect 253934 119620 253940 119632
rect 253992 119620 253998 119672
rect 254486 119620 254492 119672
rect 254544 119660 254550 119672
rect 289909 119663 289967 119669
rect 289909 119660 289921 119663
rect 254544 119632 289921 119660
rect 254544 119620 254550 119632
rect 289909 119629 289921 119632
rect 289955 119629 289967 119663
rect 289909 119623 289967 119629
rect 291841 119663 291899 119669
rect 291841 119629 291853 119663
rect 291887 119660 291899 119663
rect 291887 119632 307800 119660
rect 291887 119629 291899 119632
rect 291841 119623 291899 119629
rect 239122 119592 239128 119604
rect 61212 119564 239128 119592
rect 34974 119456 34980 119468
rect 34935 119428 34980 119456
rect 34974 119416 34980 119428
rect 35032 119416 35038 119468
rect 35158 119456 35164 119468
rect 35119 119428 35164 119456
rect 35158 119416 35164 119428
rect 35216 119416 35222 119468
rect 35342 119456 35348 119468
rect 35304 119428 35348 119456
rect 35342 119416 35348 119428
rect 35400 119416 35406 119468
rect 35529 119459 35587 119465
rect 35529 119425 35541 119459
rect 35575 119456 35587 119459
rect 35713 119459 35771 119465
rect 35713 119456 35725 119459
rect 35575 119428 35725 119456
rect 35575 119425 35587 119428
rect 35529 119419 35587 119425
rect 35713 119425 35725 119428
rect 35759 119425 35771 119459
rect 38746 119456 38752 119468
rect 38707 119428 38752 119456
rect 35713 119419 35771 119425
rect 38746 119416 38752 119428
rect 38804 119416 38810 119468
rect 61212 119465 61240 119564
rect 239122 119552 239128 119564
rect 239180 119552 239186 119604
rect 239306 119552 239312 119604
rect 239364 119592 239370 119604
rect 290550 119592 290556 119604
rect 239364 119564 290556 119592
rect 239364 119552 239370 119564
rect 290550 119552 290556 119564
rect 290608 119552 290614 119604
rect 290734 119552 290740 119604
rect 290792 119592 290798 119604
rect 307662 119592 307668 119604
rect 290792 119564 307668 119592
rect 290792 119552 290798 119564
rect 307662 119552 307668 119564
rect 307720 119552 307726 119604
rect 307772 119592 307800 119632
rect 308306 119620 308312 119672
rect 308364 119660 308370 119672
rect 314194 119660 314200 119672
rect 308364 119632 314200 119660
rect 308364 119620 308370 119632
rect 314194 119620 314200 119632
rect 314252 119620 314258 119672
rect 310422 119592 310428 119604
rect 307772 119564 310428 119592
rect 310422 119552 310428 119564
rect 310480 119552 310486 119604
rect 63494 119484 63500 119536
rect 63552 119524 63558 119536
rect 162152 119527 162210 119533
rect 63552 119496 64874 119524
rect 63552 119484 63558 119496
rect 61197 119459 61255 119465
rect 61197 119425 61209 119459
rect 61243 119425 61255 119459
rect 63678 119456 63684 119468
rect 63639 119428 63684 119456
rect 61197 119419 61255 119425
rect 63678 119416 63684 119428
rect 63736 119416 63742 119468
rect 63880 119465 63908 119496
rect 63865 119459 63923 119465
rect 63865 119425 63877 119459
rect 63911 119425 63923 119459
rect 64046 119456 64052 119468
rect 64007 119428 64052 119456
rect 63865 119419 63923 119425
rect 64046 119416 64052 119428
rect 64104 119416 64110 119468
rect 64846 119456 64874 119496
rect 142126 119496 161474 119524
rect 142126 119456 142154 119496
rect 64846 119428 142154 119456
rect 145285 119459 145343 119465
rect 145285 119425 145297 119459
rect 145331 119456 145343 119459
rect 145469 119459 145527 119465
rect 145469 119456 145481 119459
rect 145331 119428 145481 119456
rect 145331 119425 145343 119428
rect 145285 119419 145343 119425
rect 145469 119425 145481 119428
rect 145515 119425 145527 119459
rect 145650 119456 145656 119468
rect 145611 119428 145656 119456
rect 145469 119419 145527 119425
rect 145650 119416 145656 119428
rect 145708 119416 145714 119468
rect 161446 119456 161474 119496
rect 162152 119493 162164 119527
rect 162198 119524 162210 119527
rect 162198 119496 239076 119524
rect 162198 119493 162210 119496
rect 162152 119487 162210 119493
rect 215570 119456 215576 119468
rect 161446 119428 214604 119456
rect 215531 119428 215576 119456
rect 35253 119391 35311 119397
rect 35253 119357 35265 119391
rect 35299 119388 35311 119391
rect 156601 119391 156659 119397
rect 156601 119388 156613 119391
rect 35299 119360 156613 119388
rect 35299 119357 35311 119360
rect 35253 119351 35311 119357
rect 156601 119357 156613 119360
rect 156647 119357 156659 119391
rect 162394 119388 162400 119400
rect 162355 119360 162400 119388
rect 156601 119351 156659 119357
rect 162394 119348 162400 119360
rect 162452 119348 162458 119400
rect 166261 119391 166319 119397
rect 166261 119357 166273 119391
rect 166307 119388 166319 119391
rect 214469 119391 214527 119397
rect 214469 119388 214481 119391
rect 166307 119360 214481 119388
rect 166307 119357 166319 119360
rect 166261 119351 166319 119357
rect 214469 119357 214481 119360
rect 214515 119357 214527 119391
rect 214576 119388 214604 119428
rect 215570 119416 215576 119428
rect 215628 119416 215634 119468
rect 215754 119456 215760 119468
rect 215715 119428 215760 119456
rect 215754 119416 215760 119428
rect 215812 119416 215818 119468
rect 215846 119416 215852 119468
rect 215904 119456 215910 119468
rect 216122 119456 216128 119468
rect 215904 119428 215949 119456
rect 216083 119428 216128 119456
rect 215904 119416 215910 119428
rect 216122 119416 216128 119428
rect 216180 119416 216186 119468
rect 233881 119459 233939 119465
rect 233881 119456 233893 119459
rect 216232 119428 233893 119456
rect 216030 119388 216036 119400
rect 214576 119360 215800 119388
rect 215991 119360 216036 119388
rect 214469 119351 214527 119357
rect 75549 119323 75607 119329
rect 75549 119289 75561 119323
rect 75595 119320 75607 119323
rect 75733 119323 75791 119329
rect 75733 119320 75745 119323
rect 75595 119292 75745 119320
rect 75595 119289 75607 119292
rect 75549 119283 75607 119289
rect 75733 119289 75745 119292
rect 75779 119289 75791 119323
rect 75733 119283 75791 119289
rect 80977 119323 81035 119329
rect 80977 119289 80989 119323
rect 81023 119320 81035 119323
rect 81345 119323 81403 119329
rect 81345 119320 81357 119323
rect 81023 119292 81357 119320
rect 81023 119289 81035 119292
rect 80977 119283 81035 119289
rect 81345 119289 81357 119292
rect 81391 119289 81403 119323
rect 145742 119320 145748 119332
rect 145703 119292 145748 119320
rect 81345 119283 81403 119289
rect 145742 119280 145748 119292
rect 145800 119280 145806 119332
rect 215772 119320 215800 119360
rect 216030 119348 216036 119360
rect 216088 119348 216094 119400
rect 216232 119320 216260 119428
rect 233881 119425 233893 119428
rect 233927 119425 233939 119459
rect 238754 119456 238760 119468
rect 238715 119428 238760 119456
rect 233881 119419 233939 119425
rect 238754 119416 238760 119428
rect 238812 119416 238818 119468
rect 238846 119416 238852 119468
rect 238904 119456 238910 119468
rect 239048 119456 239076 119496
rect 239398 119484 239404 119536
rect 239456 119524 239462 119536
rect 253109 119527 253167 119533
rect 253109 119524 253121 119527
rect 239456 119496 253121 119524
rect 239456 119484 239462 119496
rect 253109 119493 253121 119496
rect 253155 119493 253167 119527
rect 289906 119524 289912 119536
rect 253109 119487 253167 119493
rect 253216 119496 289912 119524
rect 253216 119456 253244 119496
rect 289906 119484 289912 119496
rect 289964 119484 289970 119536
rect 290458 119524 290464 119536
rect 290292 119496 290464 119524
rect 254210 119456 254216 119468
rect 238904 119428 238949 119456
rect 239048 119428 253244 119456
rect 254171 119428 254216 119456
rect 238904 119416 238910 119428
rect 254210 119416 254216 119428
rect 254268 119416 254274 119468
rect 254305 119459 254363 119465
rect 254305 119425 254317 119459
rect 254351 119456 254363 119459
rect 255225 119459 255283 119465
rect 255225 119456 255237 119459
rect 254351 119428 255237 119456
rect 254351 119425 254363 119428
rect 254305 119419 254363 119425
rect 255225 119425 255237 119428
rect 255271 119425 255283 119459
rect 255225 119419 255283 119425
rect 258721 119459 258779 119465
rect 258721 119425 258733 119459
rect 258767 119456 258779 119459
rect 289722 119456 289728 119468
rect 258767 119428 289728 119456
rect 258767 119425 258779 119428
rect 258721 119419 258779 119425
rect 289722 119416 289728 119428
rect 289780 119416 289786 119468
rect 290292 119465 290320 119496
rect 290458 119484 290464 119496
rect 290516 119484 290522 119536
rect 291933 119527 291991 119533
rect 291933 119524 291945 119527
rect 290568 119496 291945 119524
rect 290568 119465 290596 119496
rect 291933 119493 291945 119496
rect 291979 119493 291991 119527
rect 434714 119524 434720 119536
rect 291933 119487 291991 119493
rect 292040 119496 434720 119524
rect 290277 119459 290335 119465
rect 290277 119425 290289 119459
rect 290323 119425 290335 119459
rect 290277 119419 290335 119425
rect 290553 119459 290611 119465
rect 290553 119425 290565 119459
rect 290599 119425 290611 119459
rect 290553 119419 290611 119425
rect 233329 119391 233387 119397
rect 233329 119388 233341 119391
rect 219406 119360 233341 119388
rect 151786 119292 161474 119320
rect 5902 119212 5908 119264
rect 5960 119252 5966 119264
rect 33505 119255 33563 119261
rect 33505 119252 33517 119255
rect 5960 119224 33517 119252
rect 5960 119212 5966 119224
rect 33505 119221 33517 119224
rect 33551 119221 33563 119255
rect 34882 119252 34888 119264
rect 34843 119224 34888 119252
rect 33505 119215 33563 119221
rect 34882 119212 34888 119224
rect 34940 119212 34946 119264
rect 38838 119252 38844 119264
rect 38799 119224 38844 119252
rect 38838 119212 38844 119224
rect 38896 119212 38902 119264
rect 102689 119255 102747 119261
rect 102689 119221 102701 119255
rect 102735 119252 102747 119255
rect 151786 119252 151814 119292
rect 161014 119252 161020 119264
rect 102735 119224 151814 119252
rect 160975 119224 161020 119252
rect 102735 119221 102747 119224
rect 102689 119215 102747 119221
rect 161014 119212 161020 119224
rect 161072 119212 161078 119264
rect 161446 119252 161474 119292
rect 171106 119292 180794 119320
rect 171106 119252 171134 119292
rect 172698 119252 172704 119264
rect 161446 119224 171134 119252
rect 172659 119224 172704 119252
rect 172698 119212 172704 119224
rect 172756 119212 172762 119264
rect 180766 119252 180794 119292
rect 200086 119292 215708 119320
rect 215772 119292 216260 119320
rect 216309 119323 216367 119329
rect 200086 119252 200114 119292
rect 180766 119224 200114 119252
rect 215680 119252 215708 119292
rect 216309 119289 216321 119323
rect 216355 119320 216367 119323
rect 219406 119320 219434 119360
rect 233329 119357 233341 119360
rect 233375 119357 233387 119391
rect 233329 119351 233387 119357
rect 234065 119391 234123 119397
rect 234065 119357 234077 119391
rect 234111 119388 234123 119391
rect 239030 119388 239036 119400
rect 234111 119360 239036 119388
rect 234111 119357 234123 119360
rect 234065 119351 234123 119357
rect 239030 119348 239036 119360
rect 239088 119348 239094 119400
rect 239125 119391 239183 119397
rect 239125 119357 239137 119391
rect 239171 119388 239183 119391
rect 239217 119391 239275 119397
rect 239217 119388 239229 119391
rect 239171 119360 239229 119388
rect 239171 119357 239183 119360
rect 239125 119351 239183 119357
rect 239217 119357 239229 119360
rect 239263 119357 239275 119391
rect 239217 119351 239275 119357
rect 239306 119348 239312 119400
rect 239364 119388 239370 119400
rect 239493 119391 239551 119397
rect 239364 119360 239444 119388
rect 239364 119348 239370 119360
rect 238297 119323 238355 119329
rect 238297 119320 238309 119323
rect 216355 119292 219434 119320
rect 229066 119292 238309 119320
rect 216355 119289 216367 119292
rect 216309 119283 216367 119289
rect 229066 119252 229094 119292
rect 238297 119289 238309 119292
rect 238343 119289 238355 119323
rect 239416 119320 239444 119360
rect 239493 119357 239505 119391
rect 239539 119388 239551 119391
rect 248417 119391 248475 119397
rect 248417 119388 248429 119391
rect 239539 119360 248429 119388
rect 239539 119357 239551 119360
rect 239493 119351 239551 119357
rect 248417 119357 248429 119360
rect 248463 119357 248475 119391
rect 248417 119351 248475 119357
rect 248506 119348 248512 119400
rect 248564 119388 248570 119400
rect 289817 119391 289875 119397
rect 248564 119360 277394 119388
rect 248564 119348 248570 119360
rect 253109 119323 253167 119329
rect 238297 119283 238355 119289
rect 238496 119292 239352 119320
rect 239416 119292 253060 119320
rect 215680 119224 229094 119252
rect 233329 119255 233387 119261
rect 233329 119221 233341 119255
rect 233375 119252 233387 119255
rect 238496 119252 238524 119292
rect 233375 119224 238524 119252
rect 238573 119255 238631 119261
rect 233375 119221 233387 119224
rect 233329 119215 233387 119221
rect 238573 119221 238585 119255
rect 238619 119252 238631 119255
rect 238938 119252 238944 119264
rect 238619 119224 238944 119252
rect 238619 119221 238631 119224
rect 238573 119215 238631 119221
rect 238938 119212 238944 119224
rect 238996 119212 239002 119264
rect 239033 119255 239091 119261
rect 239033 119221 239045 119255
rect 239079 119252 239091 119255
rect 239324 119252 239352 119292
rect 248230 119252 248236 119264
rect 239079 119224 239260 119252
rect 239324 119224 248236 119252
rect 239079 119221 239091 119224
rect 239033 119215 239091 119221
rect 239232 119184 239260 119224
rect 248230 119212 248236 119224
rect 248288 119212 248294 119264
rect 248325 119255 248383 119261
rect 248325 119221 248337 119255
rect 248371 119252 248383 119255
rect 253032 119252 253060 119292
rect 253109 119289 253121 119323
rect 253155 119320 253167 119323
rect 258629 119323 258687 119329
rect 258629 119320 258641 119323
rect 253155 119292 258641 119320
rect 253155 119289 253167 119292
rect 253109 119283 253167 119289
rect 258629 119289 258641 119292
rect 258675 119289 258687 119323
rect 277366 119320 277394 119360
rect 289817 119357 289829 119391
rect 289863 119388 289875 119391
rect 290185 119391 290243 119397
rect 290185 119388 290197 119391
rect 289863 119360 290197 119388
rect 289863 119357 289875 119360
rect 289817 119351 289875 119357
rect 290185 119357 290197 119360
rect 290231 119357 290243 119391
rect 290185 119351 290243 119357
rect 290366 119348 290372 119400
rect 290424 119388 290430 119400
rect 292040 119388 292068 119496
rect 434714 119484 434720 119496
rect 434772 119484 434778 119536
rect 385770 119456 385776 119468
rect 296686 119428 385776 119456
rect 290424 119360 292068 119388
rect 290424 119348 290430 119360
rect 292114 119348 292120 119400
rect 292172 119388 292178 119400
rect 296686 119388 296714 119428
rect 385770 119416 385776 119428
rect 385828 119416 385834 119468
rect 355502 119388 355508 119400
rect 292172 119360 296714 119388
rect 301516 119360 355508 119388
rect 292172 119348 292178 119360
rect 301516 119320 301544 119360
rect 355502 119348 355508 119360
rect 355560 119348 355566 119400
rect 277366 119292 301544 119320
rect 301593 119323 301651 119329
rect 258629 119283 258687 119289
rect 301593 119289 301605 119323
rect 301639 119320 301651 119323
rect 307665 119323 307723 119329
rect 307665 119320 307677 119323
rect 301639 119292 307677 119320
rect 301639 119289 301651 119292
rect 301593 119283 301651 119289
rect 307665 119289 307677 119292
rect 307711 119289 307723 119323
rect 307665 119283 307723 119289
rect 308033 119323 308091 119329
rect 308033 119289 308045 119323
rect 308079 119320 308091 119323
rect 351914 119320 351920 119332
rect 308079 119292 351920 119320
rect 308079 119289 308091 119292
rect 308033 119283 308091 119289
rect 351914 119280 351920 119292
rect 351972 119280 351978 119332
rect 258721 119255 258779 119261
rect 258721 119252 258733 119255
rect 248371 119224 252968 119252
rect 253032 119224 258733 119252
rect 248371 119221 248383 119224
rect 248325 119215 248383 119221
rect 239309 119187 239367 119193
rect 239309 119184 239321 119187
rect 239232 119156 239321 119184
rect 239309 119153 239321 119156
rect 239355 119184 239367 119187
rect 239585 119187 239643 119193
rect 239585 119184 239597 119187
rect 239355 119156 239597 119184
rect 239355 119153 239367 119156
rect 239309 119147 239367 119153
rect 239585 119153 239597 119156
rect 239631 119153 239643 119187
rect 252940 119184 252968 119224
rect 258721 119221 258733 119224
rect 258767 119221 258779 119255
rect 496538 119252 496544 119264
rect 258721 119215 258779 119221
rect 258828 119224 496544 119252
rect 253937 119187 253995 119193
rect 253937 119184 253949 119187
rect 252940 119156 253949 119184
rect 239585 119147 239643 119153
rect 253937 119153 253949 119156
rect 253983 119153 253995 119187
rect 253937 119147 253995 119153
rect 254489 119119 254547 119125
rect 254489 119085 254501 119119
rect 254535 119116 254547 119119
rect 258828 119116 258856 119224
rect 496538 119212 496544 119224
rect 496596 119212 496602 119264
rect 340966 119184 340972 119196
rect 263566 119156 289676 119184
rect 254535 119088 258856 119116
rect 258905 119119 258963 119125
rect 254535 119085 254547 119088
rect 254489 119079 254547 119085
rect 258905 119085 258917 119119
rect 258951 119116 258963 119119
rect 263566 119116 263594 119156
rect 258951 119088 263594 119116
rect 258951 119085 258963 119088
rect 258905 119079 258963 119085
rect 34606 119048 34612 119060
rect 34567 119020 34612 119048
rect 34606 119008 34612 119020
rect 34664 119008 34670 119060
rect 35713 119051 35771 119057
rect 35713 119017 35725 119051
rect 35759 119048 35771 119051
rect 48130 119048 48136 119060
rect 35759 119020 48136 119048
rect 35759 119017 35771 119020
rect 35713 119011 35771 119017
rect 48130 119008 48136 119020
rect 48188 119048 48194 119060
rect 48188 119020 234614 119048
rect 48188 119008 48194 119020
rect 4890 118940 4896 118992
rect 4948 118980 4954 118992
rect 43809 118983 43867 118989
rect 43809 118980 43821 118983
rect 4948 118952 43821 118980
rect 4948 118940 4954 118952
rect 43809 118949 43821 118952
rect 43855 118949 43867 118983
rect 43809 118943 43867 118949
rect 145650 118940 145656 118992
rect 145708 118980 145714 118992
rect 157518 118980 157524 118992
rect 145708 118952 157524 118980
rect 145708 118940 145714 118952
rect 157518 118940 157524 118952
rect 157576 118980 157582 118992
rect 168098 118980 168104 118992
rect 157576 118952 168104 118980
rect 157576 118940 157582 118952
rect 168098 118940 168104 118952
rect 168156 118940 168162 118992
rect 214469 118983 214527 118989
rect 214469 118949 214481 118983
rect 214515 118980 214527 118983
rect 216309 118983 216367 118989
rect 216309 118980 216321 118983
rect 214515 118952 216321 118980
rect 214515 118949 214527 118952
rect 214469 118943 214527 118949
rect 216309 118949 216321 118952
rect 216355 118949 216367 118983
rect 234586 118980 234614 119020
rect 238754 119008 238760 119060
rect 238812 119048 238818 119060
rect 248509 119051 248567 119057
rect 248509 119048 248521 119051
rect 238812 119020 248521 119048
rect 238812 119008 238818 119020
rect 248509 119017 248521 119020
rect 248555 119017 248567 119051
rect 289648 119048 289676 119156
rect 290660 119156 306374 119184
rect 290660 119048 290688 119156
rect 290734 119076 290740 119128
rect 290792 119116 290798 119128
rect 291933 119119 291991 119125
rect 291933 119116 291945 119119
rect 290792 119088 291945 119116
rect 290792 119076 290798 119088
rect 291933 119085 291945 119088
rect 291979 119085 291991 119119
rect 291933 119079 291991 119085
rect 297913 119119 297971 119125
rect 297913 119085 297925 119119
rect 297959 119116 297971 119119
rect 301593 119119 301651 119125
rect 301593 119116 301605 119119
rect 297959 119088 301605 119116
rect 297959 119085 297971 119088
rect 297913 119079 297971 119085
rect 301593 119085 301605 119088
rect 301639 119085 301651 119119
rect 301593 119079 301651 119085
rect 306346 119048 306374 119156
rect 308140 119156 340972 119184
rect 308140 119048 308168 119156
rect 340966 119144 340972 119156
rect 341024 119144 341030 119196
rect 308217 119119 308275 119125
rect 308217 119085 308229 119119
rect 308263 119116 308275 119119
rect 313734 119116 313740 119128
rect 308263 119088 313740 119116
rect 308263 119085 308275 119088
rect 308217 119079 308275 119085
rect 313734 119076 313740 119088
rect 313792 119076 313798 119128
rect 318150 119048 318156 119060
rect 248509 119011 248567 119017
rect 248616 119020 289584 119048
rect 289648 119020 290688 119048
rect 290752 119020 298140 119048
rect 306346 119020 308168 119048
rect 311176 119020 318156 119048
rect 248616 118980 248644 119020
rect 289556 118980 289584 119020
rect 290752 118980 290780 119020
rect 298112 118980 298140 119020
rect 311176 118980 311204 119020
rect 318150 119008 318156 119020
rect 318208 119008 318214 119060
rect 317966 118980 317972 118992
rect 234586 118952 248644 118980
rect 252388 118952 289492 118980
rect 289556 118952 290780 118980
rect 290844 118952 298048 118980
rect 298112 118952 311204 118980
rect 311268 118952 317972 118980
rect 216309 118943 216367 118949
rect 35069 118915 35127 118921
rect 35069 118881 35081 118915
rect 35115 118912 35127 118915
rect 179322 118912 179328 118924
rect 35115 118884 179328 118912
rect 35115 118881 35127 118884
rect 35069 118875 35127 118881
rect 179322 118872 179328 118884
rect 179380 118912 179386 118924
rect 179380 118884 234614 118912
rect 179380 118872 179386 118884
rect 34790 118844 34796 118856
rect 34751 118816 34796 118844
rect 34790 118804 34796 118816
rect 34848 118804 34854 118856
rect 34882 118804 34888 118856
rect 34940 118844 34946 118856
rect 35158 118844 35164 118856
rect 34940 118816 34985 118844
rect 35119 118816 35164 118844
rect 34940 118804 34946 118816
rect 35158 118804 35164 118816
rect 35216 118804 35222 118856
rect 162394 118804 162400 118856
rect 162452 118844 162458 118856
rect 180886 118844 180892 118856
rect 162452 118816 180892 118844
rect 162452 118804 162458 118816
rect 180886 118804 180892 118816
rect 180944 118804 180950 118856
rect 234586 118844 234614 118884
rect 238846 118872 238852 118924
rect 238904 118912 238910 118924
rect 252388 118912 252416 118952
rect 238904 118884 252416 118912
rect 255225 118915 255283 118921
rect 238904 118872 238910 118884
rect 255225 118881 255237 118915
rect 255271 118912 255283 118915
rect 289464 118912 289492 118952
rect 290844 118912 290872 118952
rect 255271 118884 289400 118912
rect 289464 118884 290872 118912
rect 291841 118915 291899 118921
rect 255271 118881 255283 118884
rect 255225 118875 255283 118881
rect 239309 118847 239367 118853
rect 239309 118844 239321 118847
rect 234586 118816 239321 118844
rect 239309 118813 239321 118816
rect 239355 118813 239367 118847
rect 239309 118807 239367 118813
rect 248509 118847 248567 118853
rect 248509 118813 248521 118847
rect 248555 118844 248567 118847
rect 254213 118847 254271 118853
rect 248555 118816 254072 118844
rect 248555 118813 248567 118816
rect 248509 118807 248567 118813
rect 238297 118779 238355 118785
rect 238297 118745 238309 118779
rect 238343 118776 238355 118779
rect 253937 118779 253995 118785
rect 253937 118776 253949 118779
rect 238343 118748 253949 118776
rect 238343 118745 238355 118748
rect 238297 118739 238355 118745
rect 253937 118745 253949 118748
rect 253983 118745 253995 118779
rect 254044 118776 254072 118816
rect 254213 118813 254225 118847
rect 254259 118844 254271 118847
rect 289265 118847 289323 118853
rect 289265 118844 289277 118847
rect 254259 118816 289277 118844
rect 254259 118813 254271 118816
rect 254213 118807 254271 118813
rect 289265 118813 289277 118816
rect 289311 118813 289323 118847
rect 289265 118807 289323 118813
rect 258905 118779 258963 118785
rect 258905 118776 258917 118779
rect 254044 118748 258917 118776
rect 253937 118739 253995 118745
rect 258905 118745 258917 118748
rect 258951 118745 258963 118779
rect 289372 118776 289400 118884
rect 291841 118881 291853 118915
rect 291887 118912 291899 118915
rect 297913 118915 297971 118921
rect 297913 118912 297925 118915
rect 291887 118884 297925 118912
rect 291887 118881 291899 118884
rect 291841 118875 291899 118881
rect 297913 118881 297925 118884
rect 297959 118881 297971 118915
rect 298020 118912 298048 118952
rect 311268 118912 311296 118952
rect 317966 118940 317972 118952
rect 318024 118940 318030 118992
rect 298020 118884 311296 118912
rect 297913 118875 297971 118881
rect 289449 118847 289507 118853
rect 289449 118813 289461 118847
rect 289495 118844 289507 118847
rect 307665 118847 307723 118853
rect 289495 118816 307616 118844
rect 289495 118813 289507 118816
rect 289449 118807 289507 118813
rect 291841 118779 291899 118785
rect 291841 118776 291853 118779
rect 289372 118748 291853 118776
rect 258905 118739 258963 118745
rect 291841 118745 291853 118748
rect 291887 118745 291899 118779
rect 291841 118739 291899 118745
rect 291933 118779 291991 118785
rect 291933 118745 291945 118779
rect 291979 118776 291991 118779
rect 307481 118779 307539 118785
rect 307481 118776 307493 118779
rect 291979 118748 307493 118776
rect 291979 118745 291991 118748
rect 291933 118739 291991 118745
rect 307481 118745 307493 118748
rect 307527 118745 307539 118779
rect 307588 118776 307616 118816
rect 307665 118813 307677 118847
rect 307711 118844 307723 118847
rect 318610 118844 318616 118856
rect 307711 118816 318616 118844
rect 307711 118813 307723 118816
rect 307665 118807 307723 118813
rect 318610 118804 318616 118816
rect 318668 118804 318674 118856
rect 311618 118776 311624 118788
rect 307588 118748 311624 118776
rect 307481 118739 307539 118745
rect 311618 118736 311624 118748
rect 311676 118736 311682 118788
rect 145285 118711 145343 118717
rect 145285 118677 145297 118711
rect 145331 118708 145343 118711
rect 317690 118708 317696 118720
rect 145331 118680 317696 118708
rect 145331 118677 145343 118680
rect 145285 118671 145343 118677
rect 317690 118668 317696 118680
rect 317748 118668 317754 118720
rect 9674 118600 9680 118652
rect 9732 118640 9738 118652
rect 23014 118640 23020 118652
rect 9732 118612 23020 118640
rect 9732 118600 9738 118612
rect 23014 118600 23020 118612
rect 23072 118600 23078 118652
rect 56226 118600 56232 118652
rect 56284 118640 56290 118652
rect 496262 118640 496268 118652
rect 56284 118612 496268 118640
rect 56284 118600 56290 118612
rect 496262 118600 496268 118612
rect 496320 118600 496326 118652
rect 4614 118532 4620 118584
rect 4672 118572 4678 118584
rect 16758 118572 16764 118584
rect 4672 118544 16764 118572
rect 4672 118532 4678 118544
rect 16758 118532 16764 118544
rect 16816 118532 16822 118584
rect 155586 118532 155592 118584
rect 155644 118572 155650 118584
rect 496170 118572 496176 118584
rect 155644 118544 496176 118572
rect 155644 118532 155650 118544
rect 496170 118532 496176 118544
rect 496228 118532 496234 118584
rect 162210 118464 162216 118516
rect 162268 118504 162274 118516
rect 496630 118504 496636 118516
rect 162268 118476 496636 118504
rect 162268 118464 162274 118476
rect 496630 118464 496636 118476
rect 496688 118464 496694 118516
rect 3694 118396 3700 118448
rect 3752 118436 3758 118448
rect 4890 118436 4896 118448
rect 3752 118408 4896 118436
rect 3752 118396 3758 118408
rect 4890 118396 4896 118408
rect 4948 118396 4954 118448
rect 281994 118396 282000 118448
rect 282052 118436 282058 118448
rect 467834 118436 467840 118448
rect 282052 118408 467840 118436
rect 282052 118396 282058 118408
rect 467834 118396 467840 118408
rect 467892 118396 467898 118448
rect 202230 118328 202236 118380
rect 202288 118368 202294 118380
rect 496078 118368 496084 118380
rect 202288 118340 496084 118368
rect 202288 118328 202294 118340
rect 496078 118328 496084 118340
rect 496136 118328 496142 118380
rect 6270 118260 6276 118312
rect 6328 118300 6334 118312
rect 215478 118300 215484 118312
rect 6328 118272 215484 118300
rect 6328 118260 6334 118272
rect 215478 118260 215484 118272
rect 215536 118260 215542 118312
rect 222102 118260 222108 118312
rect 222160 118300 222166 118312
rect 444006 118300 444012 118312
rect 222160 118272 444012 118300
rect 222160 118260 222166 118272
rect 444006 118260 444012 118272
rect 444064 118260 444070 118312
rect 228818 118192 228824 118244
rect 228876 118232 228882 118244
rect 438302 118232 438308 118244
rect 228876 118204 438308 118232
rect 228876 118192 228882 118204
rect 438302 118192 438308 118204
rect 438360 118192 438366 118244
rect 209130 118124 209136 118176
rect 209188 118164 209194 118176
rect 412634 118164 412640 118176
rect 209188 118136 412640 118164
rect 209188 118124 209194 118136
rect 412634 118124 412640 118136
rect 412692 118124 412698 118176
rect 122190 118056 122196 118108
rect 122248 118096 122254 118108
rect 122742 118096 122748 118108
rect 122248 118068 122748 118096
rect 122248 118056 122254 118068
rect 122742 118056 122748 118068
rect 122800 118096 122806 118108
rect 316770 118096 316776 118108
rect 122800 118068 316776 118096
rect 122800 118056 122806 118068
rect 316770 118056 316776 118068
rect 316828 118056 316834 118108
rect 308490 117988 308496 118040
rect 308548 118028 308554 118040
rect 409414 118028 409420 118040
rect 308548 118000 409420 118028
rect 308548 117988 308554 118000
rect 409414 117988 409420 118000
rect 409472 117988 409478 118040
rect 10410 117920 10416 117972
rect 10468 117960 10474 117972
rect 384298 117960 384304 117972
rect 10468 117932 384304 117960
rect 10468 117920 10474 117932
rect 384298 117920 384304 117932
rect 384356 117920 384362 117972
rect 175918 117852 175924 117904
rect 175976 117892 175982 117904
rect 316862 117892 316868 117904
rect 175976 117864 316868 117892
rect 175976 117852 175982 117864
rect 316862 117852 316868 117864
rect 316920 117852 316926 117904
rect 195330 117784 195336 117836
rect 195388 117824 195394 117836
rect 316954 117824 316960 117836
rect 195388 117796 316960 117824
rect 195388 117784 195394 117796
rect 316954 117784 316960 117796
rect 317012 117784 317018 117836
rect 295150 117716 295156 117768
rect 295208 117756 295214 117768
rect 369854 117756 369860 117768
rect 295208 117728 369860 117756
rect 295208 117716 295214 117728
rect 369854 117716 369860 117728
rect 369912 117716 369918 117768
rect 6178 117648 6184 117700
rect 6236 117688 6242 117700
rect 301590 117688 301596 117700
rect 6236 117660 301596 117688
rect 6236 117648 6242 117660
rect 301590 117648 301596 117660
rect 301648 117688 301654 117700
rect 310974 117688 310980 117700
rect 301648 117660 310980 117688
rect 301648 117648 301654 117660
rect 310974 117648 310980 117660
rect 311032 117648 311038 117700
rect 70026 117580 70032 117632
rect 70084 117620 70090 117632
rect 310422 117620 310428 117632
rect 70084 117592 310428 117620
rect 70084 117580 70090 117592
rect 310422 117580 310428 117592
rect 310480 117580 310486 117632
rect 22094 117308 22100 117360
rect 22152 117348 22158 117360
rect 23014 117348 23020 117360
rect 22152 117320 23020 117348
rect 22152 117308 22158 117320
rect 23014 117308 23020 117320
rect 23072 117308 23078 117360
rect 89254 117308 89260 117360
rect 89312 117348 89318 117360
rect 106458 117348 106464 117360
rect 89312 117320 106464 117348
rect 89312 117308 89318 117320
rect 106458 117308 106464 117320
rect 106516 117308 106522 117360
rect 451366 117280 451372 117292
rect 451424 117289 451430 117292
rect 451336 117252 451372 117280
rect 451366 117240 451372 117252
rect 451424 117243 451436 117289
rect 451642 117280 451648 117292
rect 451603 117252 451648 117280
rect 451424 117240 451430 117243
rect 451642 117240 451648 117252
rect 451700 117240 451706 117292
rect 431926 117116 450400 117144
rect 314102 117036 314108 117088
rect 314160 117076 314166 117088
rect 431926 117076 431954 117116
rect 450262 117076 450268 117088
rect 314160 117048 431954 117076
rect 450223 117048 450268 117076
rect 314160 117036 314166 117048
rect 450262 117036 450268 117048
rect 450320 117036 450326 117088
rect 450372 117076 450400 117116
rect 485225 117079 485283 117085
rect 485225 117076 485237 117079
rect 450372 117048 485237 117076
rect 485225 117045 485237 117048
rect 485271 117045 485283 117079
rect 485225 117039 485283 117045
rect 224313 116671 224371 116677
rect 224313 116637 224325 116671
rect 224359 116668 224371 116671
rect 314562 116668 314568 116680
rect 224359 116640 314568 116668
rect 224359 116637 224371 116640
rect 224313 116631 224371 116637
rect 314562 116628 314568 116640
rect 314620 116628 314626 116680
rect 209498 116560 209504 116612
rect 209556 116600 209562 116612
rect 310790 116600 310796 116612
rect 209556 116572 310796 116600
rect 209556 116560 209562 116572
rect 310790 116560 310796 116572
rect 310848 116560 310854 116612
rect 451642 116560 451648 116612
rect 451700 116600 451706 116612
rect 458174 116600 458180 116612
rect 451700 116572 458180 116600
rect 451700 116560 451706 116572
rect 458174 116560 458180 116572
rect 458232 116600 458238 116612
rect 495434 116600 495440 116612
rect 458232 116572 495440 116600
rect 458232 116560 458238 116572
rect 495434 116560 495440 116572
rect 495492 116560 495498 116612
rect 209498 115784 209504 115796
rect 209459 115756 209504 115784
rect 209498 115744 209504 115756
rect 209556 115744 209562 115796
rect 209866 115648 209872 115660
rect 209827 115620 209872 115648
rect 209866 115608 209872 115620
rect 209924 115608 209930 115660
rect 209682 115580 209688 115592
rect 209595 115552 209688 115580
rect 209682 115540 209688 115552
rect 209740 115580 209746 115592
rect 328546 115580 328552 115592
rect 209740 115552 328552 115580
rect 209740 115540 209746 115552
rect 328546 115540 328552 115552
rect 328604 115540 328610 115592
rect 315390 114860 315396 114912
rect 315448 114900 315454 114912
rect 440329 114903 440387 114909
rect 440329 114900 440341 114903
rect 315448 114872 440341 114900
rect 315448 114860 315454 114872
rect 440329 114869 440341 114872
rect 440375 114869 440387 114903
rect 440329 114863 440387 114869
rect 32585 114019 32643 114025
rect 32585 113985 32597 114019
rect 32631 114016 32643 114019
rect 89254 114016 89260 114028
rect 32631 113988 89260 114016
rect 32631 113985 32643 113988
rect 32585 113979 32643 113985
rect 89254 113976 89260 113988
rect 89312 113976 89318 114028
rect 32490 113880 32496 113892
rect 32451 113852 32496 113880
rect 32490 113840 32496 113852
rect 32548 113840 32554 113892
rect 69216 113444 74534 113472
rect 69216 113413 69244 113444
rect 69201 113407 69259 113413
rect 69201 113373 69213 113407
rect 69247 113373 69259 113407
rect 69382 113404 69388 113416
rect 69343 113376 69388 113404
rect 69201 113367 69259 113373
rect 69382 113364 69388 113376
rect 69440 113364 69446 113416
rect 74506 113404 74534 113444
rect 310238 113404 310244 113416
rect 74506 113376 310244 113404
rect 310238 113364 310244 113376
rect 310296 113364 310302 113416
rect 69017 113271 69075 113277
rect 69017 113237 69029 113271
rect 69063 113268 69075 113271
rect 346762 113268 346768 113280
rect 69063 113240 346768 113268
rect 69063 113237 69075 113240
rect 69017 113231 69075 113237
rect 346762 113228 346768 113240
rect 346820 113228 346826 113280
rect 273254 112956 273260 113008
rect 273312 112996 273318 113008
rect 405734 112996 405740 113008
rect 273312 112968 405740 112996
rect 273312 112956 273318 112968
rect 405734 112956 405740 112968
rect 405792 112956 405798 113008
rect 260282 112888 260288 112940
rect 260340 112928 260346 112940
rect 460198 112928 460204 112940
rect 260340 112900 460204 112928
rect 260340 112888 260346 112900
rect 460198 112888 460204 112900
rect 460256 112888 460262 112940
rect 266906 112820 266912 112872
rect 266964 112860 266970 112872
rect 405826 112860 405832 112872
rect 266964 112832 405832 112860
rect 266964 112820 266970 112832
rect 405826 112820 405832 112832
rect 405884 112820 405890 112872
rect 121178 112752 121184 112804
rect 121236 112792 121242 112804
rect 396718 112792 396724 112804
rect 121236 112764 396724 112792
rect 121236 112752 121242 112764
rect 396718 112752 396724 112764
rect 396776 112752 396782 112804
rect 127802 112684 127808 112736
rect 127860 112724 127866 112736
rect 418706 112724 418712 112736
rect 127860 112696 418712 112724
rect 127860 112684 127866 112696
rect 418706 112684 418712 112696
rect 418764 112684 418770 112736
rect 28442 112548 28448 112600
rect 28500 112588 28506 112600
rect 319438 112588 319444 112600
rect 28500 112560 319444 112588
rect 28500 112548 28506 112560
rect 319438 112548 319444 112560
rect 319496 112548 319502 112600
rect 81434 112480 81440 112532
rect 81492 112520 81498 112532
rect 403342 112520 403348 112532
rect 81492 112492 403348 112520
rect 81492 112480 81498 112492
rect 403342 112480 403348 112492
rect 403400 112480 403406 112532
rect 48314 112412 48320 112464
rect 48372 112452 48378 112464
rect 380158 112452 380164 112464
rect 48372 112424 380164 112452
rect 48372 112412 48378 112424
rect 380158 112412 380164 112424
rect 380216 112412 380222 112464
rect 15194 112344 15200 112396
rect 15252 112384 15258 112396
rect 370498 112384 370504 112396
rect 15252 112356 370504 112384
rect 15252 112344 15258 112356
rect 370498 112344 370504 112356
rect 370556 112344 370562 112396
rect 316678 112276 316684 112328
rect 316736 112316 316742 112328
rect 327350 112316 327356 112328
rect 316736 112288 327356 112316
rect 316736 112276 316742 112288
rect 327350 112276 327356 112288
rect 327408 112276 327414 112328
rect 328546 112248 328552 112260
rect 316006 112220 328408 112248
rect 328507 112220 328552 112248
rect 293402 112140 293408 112192
rect 293460 112180 293466 112192
rect 316006 112180 316034 112220
rect 328270 112180 328276 112192
rect 293460 112152 316034 112180
rect 325666 112152 328040 112180
rect 328231 112152 328276 112180
rect 293460 112140 293466 112152
rect 220538 111936 220544 111988
rect 220596 111976 220602 111988
rect 325666 111976 325694 112152
rect 327902 112044 327908 112056
rect 327828 112016 327908 112044
rect 220596 111948 325694 111976
rect 327721 111979 327779 111985
rect 220596 111936 220602 111948
rect 327721 111945 327733 111979
rect 327767 111976 327779 111979
rect 327828 111976 327856 112016
rect 327902 112004 327908 112016
rect 327960 112004 327966 112056
rect 327767 111948 327856 111976
rect 328012 111976 328040 112152
rect 328270 112140 328276 112152
rect 328328 112140 328334 112192
rect 328380 112180 328408 112220
rect 328546 112208 328552 112220
rect 328604 112208 328610 112260
rect 489914 112180 489920 112192
rect 328380 112152 489920 112180
rect 489914 112140 489920 112152
rect 489972 112140 489978 112192
rect 456058 111976 456064 111988
rect 328012 111948 456064 111976
rect 327767 111945 327779 111948
rect 327721 111939 327779 111945
rect 456058 111936 456064 111948
rect 456116 111936 456122 111988
rect 114554 111868 114560 111920
rect 114612 111908 114618 111920
rect 115106 111908 115112 111920
rect 114612 111880 115112 111908
rect 114612 111868 114618 111880
rect 115106 111868 115112 111880
rect 115164 111908 115170 111920
rect 393314 111908 393320 111920
rect 115164 111880 393320 111908
rect 115164 111868 115170 111880
rect 393314 111868 393320 111880
rect 393372 111868 393378 111920
rect 327258 111840 327264 111852
rect 327219 111812 327264 111840
rect 327258 111800 327264 111812
rect 327316 111800 327322 111852
rect 327350 111800 327356 111852
rect 327408 111840 327414 111852
rect 328546 111840 328552 111852
rect 327408 111812 327453 111840
rect 327644 111812 327948 111840
rect 328507 111812 328552 111840
rect 327408 111800 327414 111812
rect 132037 111775 132095 111781
rect 132037 111741 132049 111775
rect 132083 111772 132095 111775
rect 326801 111775 326859 111781
rect 326801 111772 326813 111775
rect 132083 111744 326813 111772
rect 132083 111741 132095 111744
rect 132037 111735 132095 111741
rect 326801 111741 326813 111744
rect 326847 111741 326859 111775
rect 326801 111735 326859 111741
rect 327169 111775 327227 111781
rect 327169 111741 327181 111775
rect 327215 111772 327227 111775
rect 327644 111772 327672 111812
rect 327920 111781 327948 111812
rect 328546 111800 328552 111812
rect 328604 111800 328610 111852
rect 329561 111843 329619 111849
rect 329561 111809 329573 111843
rect 329607 111840 329619 111843
rect 329745 111843 329803 111849
rect 329745 111840 329757 111843
rect 329607 111812 329757 111840
rect 329607 111809 329619 111812
rect 329561 111803 329619 111809
rect 329745 111809 329757 111812
rect 329791 111840 329803 111843
rect 337470 111840 337476 111852
rect 329791 111812 337476 111840
rect 329791 111809 329803 111812
rect 329745 111803 329803 111809
rect 337470 111800 337476 111812
rect 337528 111800 337534 111852
rect 327215 111744 327672 111772
rect 327905 111775 327963 111781
rect 327215 111741 327227 111744
rect 327169 111735 327227 111741
rect 327905 111741 327917 111775
rect 327951 111741 327963 111775
rect 327905 111735 327963 111741
rect 327997 111775 328055 111781
rect 327997 111741 328009 111775
rect 328043 111772 328055 111775
rect 494054 111772 494060 111784
rect 328043 111744 494060 111772
rect 328043 111741 328055 111744
rect 327997 111735 328055 111741
rect 494054 111732 494060 111744
rect 494112 111732 494118 111784
rect 179049 111707 179107 111713
rect 179049 111673 179061 111707
rect 179095 111704 179107 111707
rect 183373 111707 183431 111713
rect 183373 111704 183385 111707
rect 179095 111676 183385 111704
rect 179095 111673 179107 111676
rect 179049 111667 179107 111673
rect 183373 111673 183385 111676
rect 183419 111673 183431 111707
rect 183373 111667 183431 111673
rect 183462 111664 183468 111716
rect 183520 111704 183526 111716
rect 419626 111704 419632 111716
rect 183520 111676 419632 111704
rect 183520 111664 183526 111676
rect 419626 111664 419632 111676
rect 419684 111664 419690 111716
rect 168098 111596 168104 111648
rect 168156 111636 168162 111648
rect 194502 111636 194508 111648
rect 168156 111608 194508 111636
rect 168156 111596 168162 111608
rect 194502 111596 194508 111608
rect 194560 111596 194566 111648
rect 341426 111636 341432 111648
rect 224926 111608 341432 111636
rect 9030 111528 9036 111580
rect 9088 111568 9094 111580
rect 132770 111568 132776 111580
rect 9088 111540 132776 111568
rect 9088 111528 9094 111540
rect 132770 111528 132776 111540
rect 132828 111568 132834 111580
rect 135714 111568 135720 111580
rect 132828 111540 135720 111568
rect 132828 111528 132834 111540
rect 135714 111528 135720 111540
rect 135772 111528 135778 111580
rect 214558 111528 214564 111580
rect 214616 111568 214622 111580
rect 221645 111571 221703 111577
rect 221645 111568 221657 111571
rect 214616 111540 221657 111568
rect 214616 111528 214622 111540
rect 221645 111537 221657 111540
rect 221691 111568 221703 111571
rect 224926 111568 224954 111608
rect 341426 111596 341432 111608
rect 341484 111596 341490 111648
rect 480622 111636 480628 111648
rect 480583 111608 480628 111636
rect 480622 111596 480628 111608
rect 480680 111596 480686 111648
rect 221691 111540 224954 111568
rect 221691 111537 221703 111540
rect 221645 111531 221703 111537
rect 166261 111503 166319 111509
rect 166261 111469 166273 111503
rect 166307 111500 166319 111503
rect 170493 111503 170551 111509
rect 170493 111500 170505 111503
rect 166307 111472 170505 111500
rect 166307 111469 166319 111472
rect 166261 111463 166319 111469
rect 170493 111469 170505 111472
rect 170539 111469 170551 111503
rect 170493 111463 170551 111469
rect 173805 111503 173863 111509
rect 173805 111469 173817 111503
rect 173851 111500 173863 111503
rect 178957 111503 179015 111509
rect 178957 111500 178969 111503
rect 173851 111472 178969 111500
rect 173851 111469 173863 111472
rect 173805 111463 173863 111469
rect 178957 111469 178969 111472
rect 179003 111469 179015 111503
rect 178957 111463 179015 111469
rect 187789 111503 187847 111509
rect 187789 111469 187801 111503
rect 187835 111500 187847 111503
rect 194873 111503 194931 111509
rect 194873 111500 194885 111503
rect 187835 111472 194885 111500
rect 187835 111469 187847 111472
rect 187789 111463 187847 111469
rect 194873 111469 194885 111472
rect 194919 111469 194931 111503
rect 194873 111463 194931 111469
rect 84013 111435 84071 111441
rect 84013 111401 84025 111435
rect 84059 111432 84071 111435
rect 209682 111432 209688 111444
rect 84059 111404 209688 111432
rect 84059 111401 84071 111404
rect 84013 111395 84071 111401
rect 209682 111392 209688 111404
rect 209740 111392 209746 111444
rect 222749 111435 222807 111441
rect 222749 111401 222761 111435
rect 222795 111432 222807 111435
rect 416406 111432 416412 111444
rect 222795 111404 416412 111432
rect 222795 111401 222807 111404
rect 222749 111395 222807 111401
rect 416406 111392 416412 111404
rect 416464 111392 416470 111444
rect 5626 111324 5632 111376
rect 5684 111364 5690 111376
rect 173805 111367 173863 111373
rect 173805 111364 173817 111367
rect 5684 111336 173817 111364
rect 5684 111324 5690 111336
rect 173805 111333 173817 111336
rect 173851 111333 173863 111367
rect 173805 111327 173863 111333
rect 173897 111367 173955 111373
rect 173897 111333 173909 111367
rect 173943 111364 173955 111367
rect 179049 111367 179107 111373
rect 179049 111364 179061 111367
rect 173943 111336 179061 111364
rect 173943 111333 173955 111336
rect 173897 111327 173955 111333
rect 179049 111333 179061 111336
rect 179095 111333 179107 111367
rect 179049 111327 179107 111333
rect 179141 111367 179199 111373
rect 179141 111333 179153 111367
rect 179187 111364 179199 111367
rect 181346 111364 181352 111376
rect 179187 111336 181352 111364
rect 179187 111333 179199 111336
rect 179141 111327 179199 111333
rect 181346 111324 181352 111336
rect 181404 111324 181410 111376
rect 191009 111367 191067 111373
rect 191009 111364 191021 111367
rect 181456 111336 191021 111364
rect 106458 111256 106464 111308
rect 106516 111296 106522 111308
rect 162394 111296 162400 111308
rect 106516 111268 162400 111296
rect 106516 111256 106522 111268
rect 162394 111256 162400 111268
rect 162452 111256 162458 111308
rect 168374 111256 168380 111308
rect 168432 111296 168438 111308
rect 181456 111296 181484 111336
rect 191009 111333 191021 111336
rect 191055 111333 191067 111367
rect 202509 111367 202567 111373
rect 202509 111364 202521 111367
rect 191009 111327 191067 111333
rect 191116 111336 202521 111364
rect 168432 111268 181484 111296
rect 168432 111256 168438 111268
rect 181622 111256 181628 111308
rect 181680 111296 181686 111308
rect 191116 111296 191144 111336
rect 202509 111333 202521 111336
rect 202555 111333 202567 111367
rect 202509 111327 202567 111333
rect 222378 111324 222384 111376
rect 222436 111364 222442 111376
rect 417418 111364 417424 111376
rect 222436 111336 417424 111364
rect 222436 111324 222442 111336
rect 417418 111324 417424 111336
rect 417476 111324 417482 111376
rect 367094 111296 367100 111308
rect 181680 111268 191144 111296
rect 195946 111268 367100 111296
rect 181680 111256 181686 111268
rect 6638 111188 6644 111240
rect 6696 111228 6702 111240
rect 178957 111231 179015 111237
rect 6696 111200 174124 111228
rect 6696 111188 6702 111200
rect 28629 111163 28687 111169
rect 28629 111129 28641 111163
rect 28675 111160 28687 111163
rect 174096 111160 174124 111200
rect 178957 111197 178969 111231
rect 179003 111228 179015 111231
rect 179509 111231 179567 111237
rect 179509 111228 179521 111231
rect 179003 111200 179521 111228
rect 179003 111197 179015 111200
rect 178957 111191 179015 111197
rect 179509 111197 179521 111200
rect 179555 111228 179567 111231
rect 179601 111231 179659 111237
rect 179601 111228 179613 111231
rect 179555 111200 179613 111228
rect 179555 111197 179567 111200
rect 179509 111191 179567 111197
rect 179601 111197 179613 111200
rect 179647 111197 179659 111231
rect 181993 111231 182051 111237
rect 179601 111191 179659 111197
rect 179800 111200 181944 111228
rect 179141 111163 179199 111169
rect 179141 111160 179153 111163
rect 28675 111132 174032 111160
rect 174096 111132 179153 111160
rect 28675 111129 28687 111132
rect 28629 111123 28687 111129
rect 106277 111095 106335 111101
rect 106277 111061 106289 111095
rect 106323 111092 106335 111095
rect 108301 111095 108359 111101
rect 108301 111092 108313 111095
rect 106323 111064 108313 111092
rect 106323 111061 106335 111064
rect 106277 111055 106335 111061
rect 108301 111061 108313 111064
rect 108347 111061 108359 111095
rect 108301 111055 108359 111061
rect 108393 111095 108451 111101
rect 108393 111061 108405 111095
rect 108439 111092 108451 111095
rect 173897 111095 173955 111101
rect 173897 111092 173909 111095
rect 108439 111064 173909 111092
rect 108439 111061 108451 111064
rect 108393 111055 108451 111061
rect 173897 111061 173909 111064
rect 173943 111061 173955 111095
rect 174004 111092 174032 111132
rect 179141 111129 179153 111132
rect 179187 111129 179199 111163
rect 179800 111160 179828 111200
rect 179141 111123 179199 111129
rect 179248 111132 179828 111160
rect 179969 111163 180027 111169
rect 179248 111092 179276 111132
rect 179969 111129 179981 111163
rect 180015 111160 180027 111163
rect 181806 111160 181812 111172
rect 180015 111132 181812 111160
rect 180015 111129 180027 111132
rect 179969 111123 180027 111129
rect 181806 111120 181812 111132
rect 181864 111120 181870 111172
rect 181916 111160 181944 111200
rect 181993 111197 182005 111231
rect 182039 111228 182051 111231
rect 182082 111228 182088 111240
rect 182039 111200 182088 111228
rect 182039 111197 182051 111200
rect 181993 111191 182051 111197
rect 182082 111188 182088 111200
rect 182140 111228 182146 111240
rect 182818 111228 182824 111240
rect 182140 111200 182824 111228
rect 182140 111188 182146 111200
rect 182818 111188 182824 111200
rect 182876 111188 182882 111240
rect 182913 111231 182971 111237
rect 182913 111197 182925 111231
rect 182959 111228 182971 111231
rect 183097 111231 183155 111237
rect 183097 111228 183109 111231
rect 182959 111200 183109 111228
rect 182959 111197 182971 111200
rect 182913 111191 182971 111197
rect 183097 111197 183109 111200
rect 183143 111197 183155 111231
rect 183097 111191 183155 111197
rect 190089 111231 190147 111237
rect 190089 111197 190101 111231
rect 190135 111228 190147 111231
rect 190917 111231 190975 111237
rect 190917 111228 190929 111231
rect 190135 111200 190929 111228
rect 190135 111197 190147 111200
rect 190089 111191 190147 111197
rect 190917 111197 190929 111200
rect 190963 111197 190975 111231
rect 190917 111191 190975 111197
rect 191009 111231 191067 111237
rect 191009 111197 191021 111231
rect 191055 111228 191067 111231
rect 195946 111228 195974 111268
rect 367094 111256 367100 111268
rect 367152 111256 367158 111308
rect 191055 111200 195974 111228
rect 212629 111231 212687 111237
rect 191055 111197 191067 111200
rect 191009 111191 191067 111197
rect 212629 111197 212641 111231
rect 212675 111228 212687 111231
rect 213638 111228 213644 111240
rect 212675 111200 213644 111228
rect 212675 111197 212687 111200
rect 212629 111191 212687 111197
rect 213638 111188 213644 111200
rect 213696 111228 213702 111240
rect 221918 111228 221924 111240
rect 213696 111200 221924 111228
rect 213696 111188 213702 111200
rect 221918 111188 221924 111200
rect 221976 111188 221982 111240
rect 222010 111188 222016 111240
rect 222068 111228 222074 111240
rect 222933 111231 222991 111237
rect 222933 111228 222945 111231
rect 222068 111200 222945 111228
rect 222068 111188 222074 111200
rect 222933 111197 222945 111200
rect 222979 111197 222991 111231
rect 222933 111191 222991 111197
rect 273625 111231 273683 111237
rect 273625 111197 273637 111231
rect 273671 111228 273683 111231
rect 326801 111231 326859 111237
rect 273671 111200 316034 111228
rect 273671 111197 273683 111200
rect 273625 111191 273683 111197
rect 231854 111160 231860 111172
rect 181916 111132 231860 111160
rect 231854 111120 231860 111132
rect 231912 111120 231918 111172
rect 272429 111163 272487 111169
rect 272429 111129 272441 111163
rect 272475 111160 272487 111163
rect 274085 111163 274143 111169
rect 274085 111160 274097 111163
rect 272475 111132 274097 111160
rect 272475 111129 272487 111132
rect 272429 111123 272487 111129
rect 274085 111129 274097 111132
rect 274131 111129 274143 111163
rect 274085 111123 274143 111129
rect 274177 111163 274235 111169
rect 274177 111129 274189 111163
rect 274223 111160 274235 111163
rect 310330 111160 310336 111172
rect 274223 111132 310336 111160
rect 274223 111129 274235 111132
rect 274177 111123 274235 111129
rect 310330 111120 310336 111132
rect 310388 111120 310394 111172
rect 316006 111160 316034 111200
rect 326801 111197 326813 111231
rect 326847 111228 326859 111231
rect 327997 111231 328055 111237
rect 327997 111228 328009 111231
rect 326847 111200 328009 111228
rect 326847 111197 326859 111200
rect 326801 111191 326859 111197
rect 327997 111197 328009 111200
rect 328043 111197 328055 111231
rect 327997 111191 328055 111197
rect 328733 111231 328791 111237
rect 328733 111197 328745 111231
rect 328779 111228 328791 111231
rect 329745 111231 329803 111237
rect 329745 111228 329757 111231
rect 328779 111200 329757 111228
rect 328779 111197 328791 111200
rect 328733 111191 328791 111197
rect 329745 111197 329757 111200
rect 329791 111197 329803 111231
rect 472618 111228 472624 111240
rect 329745 111191 329803 111197
rect 335326 111200 472624 111228
rect 335326 111160 335354 111200
rect 472618 111188 472624 111200
rect 472676 111188 472682 111240
rect 316006 111132 335354 111160
rect 174004 111064 179276 111092
rect 173897 111055 173955 111061
rect 179322 111052 179328 111104
rect 179380 111092 179386 111104
rect 179380 111064 179425 111092
rect 179380 111052 179386 111064
rect 179874 111052 179880 111104
rect 179932 111092 179938 111104
rect 183281 111095 183339 111101
rect 183281 111092 183293 111095
rect 179932 111064 183293 111092
rect 179932 111052 179938 111064
rect 183281 111061 183293 111064
rect 183327 111061 183339 111095
rect 183281 111055 183339 111061
rect 183373 111095 183431 111101
rect 183373 111061 183385 111095
rect 183419 111092 183431 111095
rect 316586 111092 316592 111104
rect 183419 111064 316592 111092
rect 183419 111061 183431 111064
rect 183373 111055 183431 111061
rect 316586 111052 316592 111064
rect 316644 111052 316650 111104
rect 327905 111095 327963 111101
rect 327905 111061 327917 111095
rect 327951 111092 327963 111095
rect 328273 111095 328331 111101
rect 328273 111092 328285 111095
rect 327951 111064 328285 111092
rect 327951 111061 327963 111064
rect 327905 111055 327963 111061
rect 328273 111061 328285 111064
rect 328319 111061 328331 111095
rect 328273 111055 328331 111061
rect 183186 110984 183192 111036
rect 183244 111024 183250 111036
rect 183244 110996 190224 111024
rect 183244 110984 183250 110996
rect 183094 110916 183100 110968
rect 183152 110956 183158 110968
rect 187789 110959 187847 110965
rect 187789 110956 187801 110959
rect 183152 110928 187801 110956
rect 183152 110916 183158 110928
rect 187789 110925 187801 110928
rect 187835 110925 187847 110959
rect 187789 110919 187847 110925
rect 82817 110891 82875 110897
rect 82817 110857 82829 110891
rect 82863 110888 82875 110891
rect 83093 110891 83151 110897
rect 83093 110888 83105 110891
rect 82863 110860 83105 110888
rect 82863 110857 82875 110860
rect 82817 110851 82875 110857
rect 83093 110857 83105 110860
rect 83139 110857 83151 110891
rect 83093 110851 83151 110857
rect 83461 110891 83519 110897
rect 83461 110857 83473 110891
rect 83507 110888 83519 110891
rect 190089 110891 190147 110897
rect 190089 110888 190101 110891
rect 83507 110860 190101 110888
rect 83507 110857 83519 110860
rect 83461 110851 83519 110857
rect 190089 110857 190101 110860
rect 190135 110857 190147 110891
rect 190196 110888 190224 110996
rect 194796 110996 202644 111024
rect 194796 110888 194824 110996
rect 190196 110860 194824 110888
rect 194873 110891 194931 110897
rect 190089 110851 190147 110857
rect 194873 110857 194885 110891
rect 194919 110888 194931 110891
rect 202506 110888 202512 110900
rect 194919 110860 202512 110888
rect 194919 110857 194931 110860
rect 194873 110851 194931 110857
rect 202506 110848 202512 110860
rect 202564 110848 202570 110900
rect 202616 110888 202644 110996
rect 202984 110996 214236 111024
rect 202984 110888 203012 110996
rect 202616 110860 203012 110888
rect 203058 110848 203064 110900
rect 203116 110888 203122 110900
rect 214208 110888 214236 110996
rect 222672 110996 272564 111024
rect 222672 110888 222700 110996
rect 272429 110959 272487 110965
rect 272429 110956 272441 110959
rect 203116 110860 212764 110888
rect 214208 110860 222700 110888
rect 222764 110928 272441 110956
rect 203116 110848 203122 110860
rect 5258 110780 5264 110832
rect 5316 110820 5322 110832
rect 178681 110823 178739 110829
rect 178681 110820 178693 110823
rect 5316 110792 178693 110820
rect 5316 110780 5322 110792
rect 178681 110789 178693 110792
rect 178727 110789 178739 110823
rect 178681 110783 178739 110789
rect 181073 110823 181131 110829
rect 181073 110789 181085 110823
rect 181119 110820 181131 110823
rect 212629 110823 212687 110829
rect 212629 110820 212641 110823
rect 181119 110792 212641 110820
rect 181119 110789 181131 110792
rect 181073 110783 181131 110789
rect 212629 110789 212641 110792
rect 212675 110789 212687 110823
rect 212736 110820 212764 110860
rect 222764 110820 222792 110928
rect 272429 110925 272441 110928
rect 272475 110925 272487 110959
rect 272429 110919 272487 110925
rect 272536 110888 272564 110996
rect 274174 110984 274180 111036
rect 274232 111024 274238 111036
rect 314102 111024 314108 111036
rect 274232 110996 282224 111024
rect 274232 110984 274238 110996
rect 274085 110959 274143 110965
rect 274085 110925 274097 110959
rect 274131 110956 274143 110959
rect 282089 110959 282147 110965
rect 282089 110956 282101 110959
rect 274131 110928 282101 110956
rect 274131 110925 274143 110928
rect 274085 110919 274143 110925
rect 282089 110925 282101 110928
rect 282135 110925 282147 110959
rect 282089 110919 282147 110925
rect 273438 110888 273444 110900
rect 272536 110860 273444 110888
rect 273438 110848 273444 110860
rect 273496 110848 273502 110900
rect 273533 110891 273591 110897
rect 273533 110857 273545 110891
rect 273579 110888 273591 110891
rect 274634 110888 274640 110900
rect 273579 110860 274640 110888
rect 273579 110857 273591 110860
rect 273533 110851 273591 110857
rect 274634 110848 274640 110860
rect 274692 110848 274698 110900
rect 282196 110888 282224 110996
rect 286336 110996 314108 111024
rect 286336 110888 286364 110996
rect 314102 110984 314108 110996
rect 314160 110984 314166 111036
rect 286413 110959 286471 110965
rect 286413 110925 286425 110959
rect 286459 110956 286471 110959
rect 315390 110956 315396 110968
rect 286459 110928 315396 110956
rect 286459 110925 286471 110928
rect 286413 110919 286471 110925
rect 315390 110916 315396 110928
rect 315448 110916 315454 110968
rect 282196 110860 286364 110888
rect 212736 110792 222792 110820
rect 222933 110823 222991 110829
rect 212629 110783 212687 110789
rect 222933 110789 222945 110823
rect 222979 110820 222991 110823
rect 495434 110820 495440 110832
rect 222979 110792 495440 110820
rect 222979 110789 222991 110792
rect 222933 110783 222991 110789
rect 495434 110780 495440 110792
rect 495492 110780 495498 110832
rect 28445 110755 28503 110761
rect 28445 110721 28457 110755
rect 28491 110752 28503 110755
rect 28629 110755 28687 110761
rect 28629 110752 28641 110755
rect 28491 110724 28641 110752
rect 28491 110721 28503 110724
rect 28445 110715 28503 110721
rect 28629 110721 28641 110724
rect 28675 110721 28687 110755
rect 28629 110715 28687 110721
rect 50525 110755 50583 110761
rect 50525 110721 50537 110755
rect 50571 110752 50583 110755
rect 50985 110755 51043 110761
rect 50985 110752 50997 110755
rect 50571 110724 50997 110752
rect 50571 110721 50583 110724
rect 50525 110715 50583 110721
rect 50985 110721 50997 110724
rect 51031 110721 51043 110755
rect 50985 110715 51043 110721
rect 83553 110755 83611 110761
rect 83553 110721 83565 110755
rect 83599 110752 83611 110755
rect 96890 110752 96896 110764
rect 83599 110724 84194 110752
rect 96851 110724 96896 110752
rect 83599 110721 83611 110724
rect 83553 110715 83611 110721
rect 18969 110687 19027 110693
rect 18969 110684 18981 110687
rect 6886 110656 18981 110684
rect 6886 110628 6914 110656
rect 18969 110653 18981 110656
rect 19015 110653 19027 110687
rect 18969 110647 19027 110653
rect 35158 110644 35164 110696
rect 35216 110684 35222 110696
rect 82817 110687 82875 110693
rect 82817 110684 82829 110687
rect 35216 110656 82829 110684
rect 35216 110644 35222 110656
rect 82817 110653 82829 110656
rect 82863 110653 82875 110687
rect 82817 110647 82875 110653
rect 83737 110687 83795 110693
rect 83737 110653 83749 110687
rect 83783 110684 83795 110687
rect 84013 110687 84071 110693
rect 84013 110684 84025 110687
rect 83783 110656 84025 110684
rect 83783 110653 83795 110656
rect 83737 110647 83795 110653
rect 84013 110653 84025 110656
rect 84059 110653 84071 110687
rect 84166 110684 84194 110724
rect 96890 110712 96896 110724
rect 96948 110712 96954 110764
rect 106458 110752 106464 110764
rect 106419 110724 106464 110752
rect 106458 110712 106464 110724
rect 106516 110712 106522 110764
rect 106728 110755 106786 110761
rect 106728 110721 106740 110755
rect 106774 110752 106786 110755
rect 166261 110755 166319 110761
rect 166261 110752 166273 110755
rect 106774 110724 166273 110752
rect 106774 110721 106786 110724
rect 106728 110715 106786 110721
rect 166261 110721 166273 110724
rect 166307 110721 166319 110755
rect 166261 110715 166319 110721
rect 168098 110712 168104 110764
rect 168156 110752 168162 110764
rect 168285 110755 168343 110761
rect 168156 110724 168201 110752
rect 168156 110712 168162 110724
rect 168285 110721 168297 110755
rect 168331 110750 168343 110755
rect 168374 110750 168380 110764
rect 168331 110722 168380 110750
rect 168331 110721 168343 110722
rect 168285 110715 168343 110721
rect 168374 110712 168380 110722
rect 168432 110712 168438 110764
rect 170309 110755 170367 110761
rect 170309 110721 170321 110755
rect 170355 110752 170367 110755
rect 170401 110755 170459 110761
rect 170401 110752 170413 110755
rect 170355 110724 170413 110752
rect 170355 110721 170367 110724
rect 170309 110715 170367 110721
rect 170401 110721 170413 110724
rect 170447 110721 170459 110755
rect 170401 110715 170459 110721
rect 170493 110755 170551 110761
rect 170493 110721 170505 110755
rect 170539 110752 170551 110755
rect 178589 110755 178647 110761
rect 178589 110752 178601 110755
rect 170539 110724 178601 110752
rect 170539 110721 170551 110724
rect 170493 110715 170551 110721
rect 178589 110721 178601 110724
rect 178635 110721 178647 110755
rect 178589 110715 178647 110721
rect 180610 110712 180616 110764
rect 180668 110761 180674 110764
rect 180668 110752 180680 110761
rect 182634 110752 182640 110764
rect 180668 110724 180713 110752
rect 182595 110724 182640 110752
rect 180668 110715 180680 110724
rect 180668 110712 180674 110715
rect 182634 110712 182640 110724
rect 182692 110712 182698 110764
rect 182729 110755 182787 110761
rect 182729 110721 182741 110755
rect 182775 110752 182787 110755
rect 183097 110755 183155 110761
rect 183097 110752 183109 110755
rect 182775 110724 183109 110752
rect 182775 110721 182787 110724
rect 182729 110715 182787 110721
rect 183097 110721 183109 110724
rect 183143 110721 183155 110755
rect 183097 110715 183155 110721
rect 183189 110755 183247 110761
rect 183189 110721 183201 110755
rect 183235 110752 183247 110755
rect 194318 110752 194324 110764
rect 183235 110724 194324 110752
rect 183235 110721 183247 110724
rect 183189 110715 183247 110721
rect 194318 110712 194324 110724
rect 194376 110712 194382 110764
rect 194410 110712 194416 110764
rect 194468 110752 194474 110764
rect 194594 110761 194600 110764
rect 194551 110755 194600 110761
rect 194468 110724 194513 110752
rect 194468 110712 194474 110724
rect 194551 110721 194563 110755
rect 194597 110721 194600 110755
rect 194551 110715 194600 110721
rect 194594 110712 194600 110715
rect 194652 110712 194658 110764
rect 194686 110712 194692 110764
rect 194744 110752 194750 110764
rect 214374 110752 214380 110764
rect 194744 110724 214380 110752
rect 194744 110712 194750 110724
rect 214374 110712 214380 110724
rect 214432 110712 214438 110764
rect 214466 110712 214472 110764
rect 214524 110752 214530 110764
rect 214650 110752 214656 110764
rect 214524 110724 214569 110752
rect 214611 110724 214656 110752
rect 214524 110712 214530 110724
rect 214650 110712 214656 110724
rect 214708 110712 214714 110764
rect 221737 110755 221795 110761
rect 221826 110755 221884 110761
rect 221737 110721 221749 110755
rect 221783 110727 221838 110755
rect 221783 110721 221795 110727
rect 221737 110715 221795 110721
rect 221826 110721 221838 110727
rect 221872 110721 221884 110755
rect 221826 110715 221884 110721
rect 222010 110712 222016 110764
rect 222068 110752 222074 110764
rect 222068 110724 222112 110752
rect 222068 110712 222074 110724
rect 222194 110712 222200 110764
rect 222252 110752 222258 110764
rect 222252 110724 222297 110752
rect 222252 110712 222258 110724
rect 222378 110712 222384 110764
rect 222436 110752 222442 110764
rect 222436 110724 222481 110752
rect 222436 110712 222442 110724
rect 222562 110712 222568 110764
rect 222620 110752 222626 110764
rect 418982 110752 418988 110764
rect 222620 110724 418988 110752
rect 222620 110712 222626 110724
rect 418982 110712 418988 110724
rect 419040 110712 419046 110764
rect 106277 110687 106335 110693
rect 106277 110684 106289 110687
rect 84166 110656 106289 110684
rect 84013 110647 84071 110653
rect 106277 110653 106289 110656
rect 106323 110653 106335 110687
rect 106277 110647 106335 110653
rect 108301 110687 108359 110693
rect 108301 110653 108313 110687
rect 108347 110684 108359 110687
rect 179874 110684 179880 110696
rect 108347 110656 179880 110684
rect 108347 110653 108359 110656
rect 108301 110647 108359 110653
rect 179874 110644 179880 110656
rect 179932 110644 179938 110696
rect 180886 110684 180892 110696
rect 180847 110656 180892 110684
rect 180886 110644 180892 110656
rect 180944 110644 180950 110696
rect 181254 110644 181260 110696
rect 181312 110684 181318 110696
rect 181533 110687 181591 110693
rect 181533 110684 181545 110687
rect 181312 110656 181545 110684
rect 181312 110644 181318 110656
rect 181533 110653 181545 110656
rect 181579 110653 181591 110687
rect 182082 110684 182088 110696
rect 182043 110656 182088 110684
rect 181533 110647 181591 110653
rect 182082 110644 182088 110656
rect 182140 110644 182146 110696
rect 222102 110693 222108 110696
rect 183281 110687 183339 110693
rect 183281 110653 183293 110687
rect 183327 110684 183339 110687
rect 221645 110687 221703 110693
rect 221645 110684 221657 110687
rect 183327 110656 221657 110684
rect 183327 110653 183339 110656
rect 183281 110647 183339 110653
rect 221645 110653 221657 110656
rect 221691 110653 221703 110687
rect 221645 110647 221703 110653
rect 222100 110647 222108 110693
rect 222160 110684 222166 110696
rect 224957 110687 225015 110693
rect 224957 110684 224969 110687
rect 222160 110656 222200 110684
rect 222396 110656 224969 110684
rect 222102 110644 222108 110647
rect 222160 110644 222166 110656
rect 6822 110576 6828 110628
rect 6880 110588 6914 110628
rect 50985 110619 51043 110625
rect 16546 110588 35894 110616
rect 6880 110576 6886 110588
rect 4982 110508 4988 110560
rect 5040 110548 5046 110560
rect 16546 110548 16574 110588
rect 5040 110520 16574 110548
rect 35866 110548 35894 110588
rect 45526 110588 50660 110616
rect 45526 110548 45554 110588
rect 35866 110520 45554 110548
rect 50632 110548 50660 110588
rect 50985 110585 50997 110619
rect 51031 110616 51043 110619
rect 168098 110616 168104 110628
rect 51031 110588 103514 110616
rect 51031 110585 51043 110588
rect 50985 110579 51043 110585
rect 101033 110551 101091 110557
rect 101033 110548 101045 110551
rect 50632 110520 101045 110548
rect 5040 110508 5046 110520
rect 101033 110517 101045 110520
rect 101079 110517 101091 110551
rect 103486 110548 103514 110588
rect 107764 110588 161474 110616
rect 168059 110588 168104 110616
rect 107764 110548 107792 110588
rect 103486 110520 107792 110548
rect 107841 110551 107899 110557
rect 101033 110511 101091 110517
rect 107841 110517 107853 110551
rect 107887 110548 107899 110551
rect 108393 110551 108451 110557
rect 108393 110548 108405 110551
rect 107887 110520 108405 110548
rect 107887 110517 107899 110520
rect 107841 110511 107899 110517
rect 108393 110517 108405 110520
rect 108439 110517 108451 110551
rect 108393 110511 108451 110517
rect 131485 110551 131543 110557
rect 131485 110517 131497 110551
rect 131531 110548 131543 110551
rect 132037 110551 132095 110557
rect 132037 110548 132049 110551
rect 131531 110520 132049 110548
rect 131531 110517 131543 110520
rect 131485 110511 131543 110517
rect 132037 110517 132049 110520
rect 132083 110517 132095 110551
rect 137186 110548 137192 110560
rect 137147 110520 137192 110548
rect 132037 110511 132095 110517
rect 137186 110508 137192 110520
rect 137244 110508 137250 110560
rect 161446 110548 161474 110588
rect 168098 110576 168104 110588
rect 168156 110576 168162 110628
rect 191009 110619 191067 110625
rect 168208 110588 180012 110616
rect 168208 110548 168236 110588
rect 170214 110548 170220 110560
rect 161446 110520 168236 110548
rect 170175 110520 170220 110548
rect 170214 110508 170220 110520
rect 170272 110508 170278 110560
rect 170401 110551 170459 110557
rect 170401 110517 170413 110551
rect 170447 110548 170459 110551
rect 179506 110548 179512 110560
rect 170447 110520 179368 110548
rect 179467 110520 179512 110548
rect 170447 110517 170459 110520
rect 170401 110511 170459 110517
rect 179340 110344 179368 110520
rect 179506 110508 179512 110520
rect 179564 110508 179570 110560
rect 179984 110548 180012 110588
rect 180904 110588 190960 110616
rect 180904 110548 180932 110588
rect 190454 110548 190460 110560
rect 179984 110520 180932 110548
rect 180996 110520 190224 110548
rect 190415 110520 190460 110548
rect 180996 110344 181024 110520
rect 179340 110316 181024 110344
rect 190196 110344 190224 110520
rect 190454 110508 190460 110520
rect 190512 110508 190518 110560
rect 190932 110548 190960 110588
rect 191009 110585 191021 110619
rect 191055 110616 191067 110619
rect 194597 110619 194655 110625
rect 194597 110616 194609 110619
rect 191055 110588 194609 110616
rect 191055 110585 191067 110588
rect 191009 110579 191067 110585
rect 194597 110585 194609 110588
rect 194643 110585 194655 110619
rect 222396 110616 222424 110656
rect 224957 110653 224969 110656
rect 225003 110653 225015 110687
rect 224957 110647 225015 110653
rect 225233 110687 225291 110693
rect 225233 110653 225245 110687
rect 225279 110684 225291 110687
rect 273438 110684 273444 110696
rect 225279 110656 273444 110684
rect 225279 110653 225291 110656
rect 225233 110647 225291 110653
rect 273438 110644 273444 110656
rect 273496 110644 273502 110696
rect 273622 110644 273628 110696
rect 273680 110684 273686 110696
rect 273680 110656 273725 110684
rect 273680 110644 273686 110656
rect 273806 110644 273812 110696
rect 273864 110684 273870 110696
rect 274177 110687 274235 110693
rect 274177 110684 274189 110687
rect 273864 110656 274189 110684
rect 273864 110644 273870 110656
rect 274177 110653 274189 110656
rect 274223 110653 274235 110687
rect 274177 110647 274235 110653
rect 282089 110687 282147 110693
rect 282089 110653 282101 110687
rect 282135 110684 282147 110687
rect 286413 110687 286471 110693
rect 286413 110684 286425 110687
rect 282135 110656 286425 110684
rect 282135 110653 282147 110656
rect 282089 110647 282147 110653
rect 286413 110653 286425 110656
rect 286459 110653 286471 110687
rect 286413 110647 286471 110653
rect 286505 110687 286563 110693
rect 286505 110653 286517 110687
rect 286551 110684 286563 110687
rect 409046 110684 409052 110696
rect 286551 110656 409052 110684
rect 286551 110653 286563 110656
rect 286505 110647 286563 110653
rect 409046 110644 409052 110656
rect 409104 110644 409110 110696
rect 222749 110619 222807 110625
rect 222749 110616 222761 110619
rect 194597 110579 194655 110585
rect 195946 110588 222424 110616
rect 222488 110588 222761 110616
rect 195946 110548 195974 110588
rect 202693 110551 202751 110557
rect 202693 110548 202705 110551
rect 190932 110520 195974 110548
rect 202616 110520 202705 110548
rect 202509 110483 202567 110489
rect 190564 110452 194272 110480
rect 190564 110344 190592 110452
rect 190196 110316 190592 110344
rect 194244 110344 194272 110452
rect 194796 110452 202460 110480
rect 194796 110344 194824 110452
rect 202432 110412 202460 110452
rect 202509 110449 202521 110483
rect 202555 110480 202567 110483
rect 202616 110480 202644 110520
rect 202693 110517 202705 110520
rect 202739 110517 202751 110551
rect 214374 110548 214380 110560
rect 202693 110511 202751 110517
rect 202984 110520 214380 110548
rect 202555 110452 202644 110480
rect 202555 110449 202567 110452
rect 202509 110443 202567 110449
rect 202432 110384 202552 110412
rect 194244 110316 194824 110344
rect 202524 110344 202552 110384
rect 202984 110344 203012 110520
rect 214374 110508 214380 110520
rect 214432 110508 214438 110560
rect 214466 110508 214472 110560
rect 214524 110548 214530 110560
rect 222378 110548 222384 110560
rect 214524 110520 222384 110548
rect 214524 110508 214530 110520
rect 222378 110508 222384 110520
rect 222436 110508 222442 110560
rect 222488 110557 222516 110588
rect 222749 110585 222761 110588
rect 222795 110585 222807 110619
rect 310882 110616 310888 110628
rect 222749 110579 222807 110585
rect 234586 110588 310888 110616
rect 222473 110551 222531 110557
rect 222473 110517 222485 110551
rect 222519 110517 222531 110551
rect 222473 110511 222531 110517
rect 224957 110483 225015 110489
rect 224957 110449 224969 110483
rect 225003 110480 225015 110483
rect 234586 110480 234614 110588
rect 310882 110576 310888 110588
rect 310940 110576 310946 110628
rect 273162 110548 273168 110560
rect 273123 110520 273168 110548
rect 273162 110508 273168 110520
rect 273220 110508 273226 110560
rect 286229 110551 286287 110557
rect 286229 110517 286241 110551
rect 286275 110548 286287 110551
rect 311158 110548 311164 110560
rect 286275 110520 311164 110548
rect 286275 110517 286287 110520
rect 286229 110511 286287 110517
rect 311158 110508 311164 110520
rect 311216 110508 311222 110560
rect 286505 110483 286563 110489
rect 286505 110480 286517 110483
rect 225003 110452 234614 110480
rect 274008 110452 285996 110480
rect 225003 110449 225015 110452
rect 224957 110443 225015 110449
rect 202524 110316 203012 110344
rect 273438 110304 273444 110356
rect 273496 110344 273502 110356
rect 274008 110344 274036 110452
rect 273496 110316 274036 110344
rect 285968 110344 285996 110452
rect 286336 110452 286517 110480
rect 286336 110344 286364 110452
rect 286505 110449 286517 110452
rect 286551 110449 286563 110483
rect 286505 110443 286563 110449
rect 285968 110316 286364 110344
rect 273496 110304 273502 110316
rect 178681 110279 178739 110285
rect 178681 110245 178693 110279
rect 178727 110276 178739 110279
rect 181073 110279 181131 110285
rect 181073 110276 181085 110279
rect 178727 110248 181085 110276
rect 178727 110245 178739 110248
rect 178681 110239 178739 110245
rect 181073 110245 181085 110248
rect 181119 110245 181131 110279
rect 181073 110239 181131 110245
rect 221645 110279 221703 110285
rect 221645 110245 221657 110279
rect 221691 110276 221703 110279
rect 225233 110279 225291 110285
rect 225233 110276 225245 110279
rect 221691 110248 225245 110276
rect 221691 110245 221703 110248
rect 221645 110239 221703 110245
rect 225233 110245 225245 110248
rect 225279 110245 225291 110279
rect 225233 110239 225291 110245
rect 178589 110211 178647 110217
rect 178589 110177 178601 110211
rect 178635 110208 178647 110211
rect 183189 110211 183247 110217
rect 183189 110208 183201 110211
rect 178635 110180 183201 110208
rect 178635 110177 178647 110180
rect 178589 110171 178647 110177
rect 183189 110177 183201 110180
rect 183235 110177 183247 110211
rect 183189 110171 183247 110177
rect 8570 109692 8576 109744
rect 8628 109732 8634 109744
rect 22094 109732 22100 109744
rect 8628 109704 22100 109732
rect 8628 109692 8634 109704
rect 22094 109692 22100 109704
rect 22152 109692 22158 109744
rect 8478 109284 8484 109336
rect 8536 109324 8542 109336
rect 20714 109324 20720 109336
rect 8536 109296 20720 109324
rect 8536 109284 8542 109296
rect 20714 109284 20720 109296
rect 20772 109324 20778 109336
rect 21542 109324 21548 109336
rect 20772 109296 21548 109324
rect 20772 109284 20778 109296
rect 21542 109284 21548 109296
rect 21600 109284 21606 109336
rect 180886 109324 180892 109336
rect 161446 109296 180892 109324
rect 7006 109148 7012 109200
rect 7064 109188 7070 109200
rect 8662 109188 8668 109200
rect 7064 109160 8668 109188
rect 7064 109148 7070 109160
rect 8662 109148 8668 109160
rect 8720 109148 8726 109200
rect 8662 109012 8668 109064
rect 8720 109052 8726 109064
rect 161446 109052 161474 109296
rect 180886 109284 180892 109296
rect 180944 109284 180950 109336
rect 453022 109188 453028 109200
rect 452983 109160 453028 109188
rect 453022 109148 453028 109160
rect 453080 109148 453086 109200
rect 8720 109024 161474 109052
rect 453209 109055 453267 109061
rect 8720 109012 8726 109024
rect 453209 109021 453221 109055
rect 453255 109052 453267 109055
rect 470594 109052 470600 109064
rect 453255 109024 470600 109052
rect 453255 109021 453267 109024
rect 453209 109015 453267 109021
rect 470594 109012 470600 109024
rect 470652 109012 470658 109064
rect 5074 108536 5080 108588
rect 5132 108576 5138 108588
rect 315206 108576 315212 108588
rect 5132 108548 315212 108576
rect 5132 108536 5138 108548
rect 315206 108536 315212 108548
rect 315264 108536 315270 108588
rect 8938 108468 8944 108520
rect 8996 108508 9002 108520
rect 366726 108508 366732 108520
rect 8996 108480 366732 108508
rect 8996 108468 9002 108480
rect 366726 108468 366732 108480
rect 366784 108468 366790 108520
rect 8386 108400 8392 108452
rect 8444 108440 8450 108452
rect 368014 108440 368020 108452
rect 8444 108412 368020 108440
rect 8444 108400 8450 108412
rect 368014 108400 368020 108412
rect 368072 108400 368078 108452
rect 7098 108332 7104 108384
rect 7156 108372 7162 108384
rect 491294 108372 491300 108384
rect 7156 108344 491300 108372
rect 7156 108332 7162 108344
rect 491294 108332 491300 108344
rect 491352 108332 491358 108384
rect 5166 108264 5172 108316
rect 5224 108304 5230 108316
rect 416590 108304 416596 108316
rect 5224 108276 416596 108304
rect 5224 108264 5230 108276
rect 416590 108264 416596 108276
rect 416648 108264 416654 108316
rect 317230 107924 317236 107976
rect 317288 107964 317294 107976
rect 419353 107967 419411 107973
rect 419353 107964 419365 107967
rect 317288 107936 419365 107964
rect 317288 107924 317294 107936
rect 419353 107933 419365 107936
rect 419399 107933 419411 107967
rect 419534 107964 419540 107976
rect 419495 107936 419540 107964
rect 419353 107927 419411 107933
rect 419534 107924 419540 107936
rect 419592 107924 419598 107976
rect 471882 107924 471888 107976
rect 471940 107964 471946 107976
rect 496357 107967 496415 107973
rect 496357 107964 496369 107967
rect 471940 107936 496369 107964
rect 471940 107924 471946 107936
rect 496357 107933 496369 107936
rect 496403 107933 496415 107967
rect 496357 107927 496415 107933
rect 317046 107788 317052 107840
rect 317104 107828 317110 107840
rect 419721 107831 419779 107837
rect 419721 107828 419733 107831
rect 317104 107800 419733 107828
rect 317104 107788 317110 107800
rect 419721 107797 419733 107800
rect 419767 107797 419779 107831
rect 419721 107791 419779 107797
rect 9490 107652 9496 107704
rect 9548 107692 9554 107704
rect 312722 107692 312728 107704
rect 9548 107664 312728 107692
rect 9548 107652 9554 107664
rect 312722 107652 312728 107664
rect 312780 107652 312786 107704
rect 358078 106292 358084 106344
rect 358136 106332 358142 106344
rect 456981 106335 457039 106341
rect 456981 106332 456993 106335
rect 358136 106304 456993 106332
rect 358136 106292 358142 106304
rect 456981 106301 456993 106304
rect 457027 106301 457039 106335
rect 456981 106295 457039 106301
rect 368382 105448 368388 105460
rect 368343 105420 368388 105448
rect 368382 105408 368388 105420
rect 368440 105408 368446 105460
rect 368569 105315 368627 105321
rect 368569 105281 368581 105315
rect 368615 105312 368627 105315
rect 372614 105312 372620 105324
rect 368615 105284 372620 105312
rect 368615 105281 368627 105284
rect 368569 105275 368627 105281
rect 372614 105272 372620 105284
rect 372672 105272 372678 105324
rect 317966 105068 317972 105120
rect 318024 105108 318030 105120
rect 368382 105108 368388 105120
rect 318024 105080 368388 105108
rect 318024 105068 318030 105080
rect 368382 105068 368388 105080
rect 368440 105068 368446 105120
rect 344646 102144 344652 102196
rect 344704 102184 344710 102196
rect 495526 102184 495532 102196
rect 344704 102156 495532 102184
rect 344704 102144 344710 102156
rect 495526 102144 495532 102156
rect 495584 102144 495590 102196
rect 2958 101056 2964 101108
rect 3016 101096 3022 101108
rect 3513 101099 3571 101105
rect 3513 101096 3525 101099
rect 3016 101068 3525 101096
rect 3016 101056 3022 101068
rect 3513 101065 3525 101068
rect 3559 101065 3571 101099
rect 3694 101096 3700 101108
rect 3655 101068 3700 101096
rect 3513 101059 3571 101065
rect 3694 101056 3700 101068
rect 3752 101056 3758 101108
rect 3605 101031 3663 101037
rect 3605 100997 3617 101031
rect 3651 101028 3663 101031
rect 9490 101028 9496 101040
rect 3651 101000 9496 101028
rect 3651 100997 3663 101000
rect 3605 100991 3663 100997
rect 9490 100988 9496 101000
rect 9548 100988 9554 101040
rect 3881 100827 3939 100833
rect 3881 100793 3893 100827
rect 3927 100824 3939 100827
rect 4982 100824 4988 100836
rect 3927 100796 4988 100824
rect 3927 100793 3939 100796
rect 3881 100787 3939 100793
rect 4982 100784 4988 100796
rect 5040 100784 5046 100836
rect 3326 100756 3332 100768
rect 3287 100728 3332 100756
rect 3326 100716 3332 100728
rect 3384 100716 3390 100768
rect 5258 100716 5264 100768
rect 5316 100756 5322 100768
rect 6178 100756 6184 100768
rect 5316 100728 6184 100756
rect 5316 100716 5322 100728
rect 6178 100716 6184 100728
rect 6236 100716 6242 100768
rect 388438 100716 388444 100768
rect 388496 100756 388502 100768
rect 487893 100759 487951 100765
rect 487893 100756 487905 100759
rect 388496 100728 487905 100756
rect 388496 100716 388502 100728
rect 487893 100725 487905 100728
rect 487939 100725 487951 100759
rect 487893 100719 487951 100725
rect 396626 99220 396632 99272
rect 396684 99260 396690 99272
rect 458174 99260 458180 99272
rect 396684 99232 458036 99260
rect 458135 99232 458180 99260
rect 396684 99220 396690 99232
rect 440878 99152 440884 99204
rect 440936 99192 440942 99204
rect 457910 99195 457968 99201
rect 457910 99192 457922 99195
rect 440936 99164 457922 99192
rect 440936 99152 440942 99164
rect 457910 99161 457922 99164
rect 457956 99161 457968 99195
rect 458008 99192 458036 99232
rect 458174 99220 458180 99232
rect 458232 99220 458238 99272
rect 495526 99260 495532 99272
rect 460906 99232 495532 99260
rect 460906 99192 460934 99232
rect 495526 99220 495532 99232
rect 495584 99220 495590 99272
rect 458008 99164 460934 99192
rect 457910 99155 457968 99161
rect 456794 99124 456800 99136
rect 456755 99096 456800 99124
rect 456794 99084 456800 99096
rect 456852 99084 456858 99136
rect 432598 93780 432604 93832
rect 432656 93820 432662 93832
rect 495526 93820 495532 93832
rect 432656 93792 495532 93820
rect 432656 93780 432662 93792
rect 495526 93780 495532 93792
rect 495584 93780 495590 93832
rect 436738 90108 436744 90160
rect 436796 90148 436802 90160
rect 438826 90151 438884 90157
rect 438826 90148 438838 90151
rect 436796 90120 438838 90148
rect 436796 90108 436802 90120
rect 438826 90117 438838 90120
rect 438872 90117 438884 90151
rect 438826 90111 438884 90117
rect 433978 90040 433984 90092
rect 434036 90080 434042 90092
rect 438581 90083 438639 90089
rect 438581 90080 438593 90083
rect 434036 90052 438593 90080
rect 434036 90040 434042 90052
rect 438581 90049 438593 90052
rect 438627 90049 438639 90083
rect 438581 90043 438639 90049
rect 318610 89836 318616 89888
rect 318668 89876 318674 89888
rect 439958 89876 439964 89888
rect 318668 89848 439964 89876
rect 318668 89836 318674 89848
rect 439958 89836 439964 89848
rect 440016 89836 440022 89888
rect 5350 89632 5356 89684
rect 5408 89672 5414 89684
rect 8018 89672 8024 89684
rect 5408 89644 8024 89672
rect 5408 89632 5414 89644
rect 8018 89632 8024 89644
rect 8076 89632 8082 89684
rect 348418 89632 348424 89684
rect 348476 89672 348482 89684
rect 495526 89672 495532 89684
rect 348476 89644 495532 89672
rect 348476 89632 348482 89644
rect 495526 89632 495532 89644
rect 495584 89632 495590 89684
rect 312538 85756 312544 85808
rect 312596 85796 312602 85808
rect 380897 85799 380955 85805
rect 380897 85796 380909 85799
rect 312596 85768 380909 85796
rect 312596 85756 312602 85768
rect 380897 85765 380909 85768
rect 380943 85765 380955 85799
rect 380897 85759 380955 85765
rect 382182 85756 382188 85808
rect 382240 85756 382246 85808
rect 312814 85688 312820 85740
rect 312872 85728 312878 85740
rect 382093 85731 382151 85737
rect 382093 85728 382105 85731
rect 312872 85700 382105 85728
rect 312872 85688 312878 85700
rect 382093 85697 382105 85700
rect 382139 85697 382151 85731
rect 382200 85728 382228 85756
rect 382200 85700 382320 85728
rect 382093 85691 382151 85697
rect 382292 85669 382320 85700
rect 380897 85663 380955 85669
rect 380897 85629 380909 85663
rect 380943 85660 380955 85663
rect 382185 85663 382243 85669
rect 382185 85660 382197 85663
rect 380943 85632 382197 85660
rect 380943 85629 380955 85632
rect 380897 85623 380955 85629
rect 382185 85629 382197 85632
rect 382231 85629 382243 85663
rect 382185 85623 382243 85629
rect 382277 85663 382335 85669
rect 382277 85629 382289 85663
rect 382323 85629 382335 85663
rect 382277 85623 382335 85629
rect 327718 85552 327724 85604
rect 327776 85592 327782 85604
rect 381725 85595 381783 85601
rect 381725 85592 381737 85595
rect 327776 85564 381737 85592
rect 327776 85552 327782 85564
rect 381725 85561 381737 85564
rect 381771 85561 381783 85595
rect 381725 85555 381783 85561
rect 311986 85484 311992 85536
rect 312044 85524 312050 85536
rect 312906 85524 312912 85536
rect 312044 85496 312912 85524
rect 312044 85484 312050 85496
rect 312906 85484 312912 85496
rect 312964 85484 312970 85536
rect 310149 84779 310207 84785
rect 310149 84745 310161 84779
rect 310195 84776 310207 84779
rect 318058 84776 318064 84788
rect 310195 84748 318064 84776
rect 310195 84745 310207 84748
rect 310149 84739 310207 84745
rect 318058 84736 318064 84748
rect 318116 84736 318122 84788
rect 310241 84643 310299 84649
rect 310241 84609 310253 84643
rect 310287 84640 310299 84643
rect 369118 84640 369124 84652
rect 310287 84612 369124 84640
rect 310287 84609 310299 84612
rect 310241 84603 310299 84609
rect 369118 84600 369124 84612
rect 369176 84600 369182 84652
rect 8846 79880 8852 79892
rect 8807 79852 8852 79880
rect 8846 79840 8852 79852
rect 8904 79840 8910 79892
rect 9122 79772 9128 79824
rect 9180 79812 9186 79824
rect 9180 79784 9352 79812
rect 9180 79772 9186 79784
rect 6178 79704 6184 79756
rect 6236 79744 6242 79756
rect 9217 79747 9275 79753
rect 9217 79744 9229 79747
rect 6236 79716 9229 79744
rect 6236 79704 6242 79716
rect 9217 79713 9229 79716
rect 9263 79713 9275 79747
rect 9217 79707 9275 79713
rect 8938 79676 8944 79688
rect 8899 79648 8944 79676
rect 8938 79636 8944 79648
rect 8996 79636 9002 79688
rect 9122 79676 9128 79688
rect 9083 79648 9128 79676
rect 9122 79636 9128 79648
rect 9180 79636 9186 79688
rect 9324 79685 9352 79784
rect 9310 79679 9368 79685
rect 9310 79645 9322 79679
rect 9356 79645 9368 79679
rect 9310 79639 9368 79645
rect 9493 79679 9551 79685
rect 9493 79645 9505 79679
rect 9539 79645 9551 79679
rect 9493 79639 9551 79645
rect 8294 79568 8300 79620
rect 8352 79608 8358 79620
rect 9508 79608 9536 79639
rect 8352 79580 9536 79608
rect 8352 79568 8358 79580
rect 443086 79268 443092 79280
rect 443047 79240 443092 79268
rect 443086 79228 443092 79240
rect 443144 79228 443150 79280
rect 442902 79200 442908 79212
rect 442863 79172 442908 79200
rect 442902 79160 442908 79172
rect 442960 79160 442966 79212
rect 443178 78996 443184 79008
rect 443139 78968 443184 78996
rect 443178 78956 443184 78968
rect 443236 78956 443242 79008
rect 338040 78696 338344 78724
rect 337746 78656 337752 78668
rect 337659 78628 337752 78656
rect 337746 78616 337752 78628
rect 337804 78656 337810 78668
rect 338040 78656 338068 78696
rect 338206 78656 338212 78668
rect 337804 78628 338068 78656
rect 338167 78628 338212 78656
rect 337804 78616 337810 78628
rect 338206 78616 338212 78628
rect 338264 78616 338270 78668
rect 338316 78656 338344 78696
rect 429838 78656 429844 78668
rect 338316 78628 429844 78656
rect 429838 78616 429844 78628
rect 429896 78616 429902 78668
rect 469858 78656 469864 78668
rect 469819 78628 469864 78656
rect 469858 78616 469864 78628
rect 469916 78616 469922 78668
rect 327810 78548 327816 78600
rect 327868 78588 327874 78600
rect 337657 78591 337715 78597
rect 337657 78588 337669 78591
rect 327868 78560 337669 78588
rect 327868 78548 327874 78560
rect 337657 78557 337669 78560
rect 337703 78557 337715 78591
rect 337657 78551 337715 78557
rect 337933 78591 337991 78597
rect 337933 78557 337945 78591
rect 337979 78557 337991 78591
rect 337933 78551 337991 78557
rect 337948 78520 337976 78551
rect 338022 78548 338028 78600
rect 338080 78588 338086 78600
rect 339310 78597 339316 78600
rect 339267 78591 339316 78597
rect 338080 78560 339172 78588
rect 338080 78548 338086 78560
rect 337948 78492 338896 78520
rect 338868 78461 338896 78492
rect 338853 78455 338911 78461
rect 338853 78421 338865 78455
rect 338899 78421 338911 78455
rect 339144 78452 339172 78560
rect 339267 78557 339279 78591
rect 339313 78557 339316 78591
rect 339267 78551 339316 78557
rect 339310 78548 339316 78551
rect 339368 78588 339374 78600
rect 469582 78588 469588 78600
rect 339368 78560 345014 78588
rect 469543 78560 469588 78588
rect 339368 78548 339374 78560
rect 344986 78520 345014 78560
rect 469582 78548 469588 78560
rect 469640 78548 469646 78600
rect 469674 78548 469680 78600
rect 469732 78588 469738 78600
rect 469953 78591 470011 78597
rect 469732 78560 469777 78588
rect 469732 78548 469738 78560
rect 469953 78557 469965 78591
rect 469999 78588 470011 78591
rect 473722 78588 473728 78600
rect 469999 78560 473728 78588
rect 469999 78557 470011 78560
rect 469953 78551 470011 78557
rect 473722 78548 473728 78560
rect 473780 78548 473786 78600
rect 406378 78520 406384 78532
rect 344986 78492 406384 78520
rect 406378 78480 406384 78492
rect 406436 78480 406442 78532
rect 469398 78452 469404 78464
rect 339144 78424 345014 78452
rect 469359 78424 469404 78452
rect 338853 78415 338911 78421
rect 344986 78248 345014 78424
rect 469398 78412 469404 78424
rect 469456 78412 469462 78464
rect 442534 78248 442540 78260
rect 344986 78220 442540 78248
rect 442534 78208 442540 78220
rect 442592 78208 442598 78260
rect 2774 76916 2780 76968
rect 2832 76956 2838 76968
rect 4706 76956 4712 76968
rect 2832 76928 4712 76956
rect 2832 76916 2838 76928
rect 4706 76916 4712 76928
rect 4764 76916 4770 76968
rect 429838 75528 429844 75540
rect 429799 75500 429844 75528
rect 429838 75488 429844 75500
rect 429896 75488 429902 75540
rect 429654 75324 429660 75336
rect 429615 75296 429660 75324
rect 429654 75284 429660 75296
rect 429712 75284 429718 75336
rect 362218 72632 362224 72684
rect 362276 72672 362282 72684
rect 378781 72675 378839 72681
rect 378781 72672 378793 72675
rect 362276 72644 378793 72672
rect 362276 72632 362282 72644
rect 378781 72641 378793 72644
rect 378827 72641 378839 72675
rect 378781 72635 378839 72641
rect 370498 72564 370504 72616
rect 370556 72604 370562 72616
rect 378873 72607 378931 72613
rect 378873 72604 378885 72607
rect 370556 72576 378885 72604
rect 370556 72564 370562 72576
rect 378873 72573 378885 72576
rect 378919 72573 378931 72607
rect 378873 72567 378931 72573
rect 378962 72564 378968 72616
rect 379020 72604 379026 72616
rect 379020 72576 379065 72604
rect 379020 72564 379026 72576
rect 367462 72428 367468 72480
rect 367520 72468 367526 72480
rect 378413 72471 378471 72477
rect 378413 72468 378425 72471
rect 367520 72440 378425 72468
rect 367520 72428 367526 72440
rect 378413 72437 378425 72440
rect 378459 72437 378471 72471
rect 378413 72431 378471 72437
rect 378962 72428 378968 72480
rect 379020 72468 379026 72480
rect 382182 72468 382188 72480
rect 379020 72440 382188 72468
rect 379020 72428 379026 72440
rect 382182 72428 382188 72440
rect 382240 72468 382246 72480
rect 418430 72468 418436 72480
rect 382240 72440 418436 72468
rect 382240 72428 382246 72440
rect 418430 72428 418436 72440
rect 418488 72428 418494 72480
rect 496446 72264 496452 72276
rect 496407 72236 496452 72264
rect 496446 72224 496452 72236
rect 496504 72224 496510 72276
rect 359458 70388 359464 70440
rect 359516 70428 359522 70440
rect 394145 70431 394203 70437
rect 394145 70428 394157 70431
rect 359516 70400 394157 70428
rect 359516 70388 359522 70400
rect 394145 70397 394157 70400
rect 394191 70397 394203 70431
rect 394145 70391 394203 70397
rect 376202 67532 376208 67584
rect 376260 67572 376266 67584
rect 376662 67572 376668 67584
rect 376260 67544 376668 67572
rect 376260 67532 376266 67544
rect 376662 67532 376668 67544
rect 376720 67572 376726 67584
rect 429654 67572 429660 67584
rect 376720 67544 429660 67572
rect 376720 67532 376726 67544
rect 429654 67532 429660 67544
rect 429712 67532 429718 67584
rect 310054 67328 310060 67380
rect 310112 67368 310118 67380
rect 310112 67340 310157 67368
rect 310112 67328 310118 67340
rect 310241 67235 310299 67241
rect 310241 67201 310253 67235
rect 310287 67232 310299 67235
rect 339310 67232 339316 67244
rect 310287 67204 339316 67232
rect 310287 67201 310299 67204
rect 310241 67195 310299 67201
rect 339310 67192 339316 67204
rect 339368 67192 339374 67244
rect 314102 66580 314108 66632
rect 314160 66620 314166 66632
rect 360289 66623 360347 66629
rect 360289 66620 360301 66623
rect 314160 66592 360301 66620
rect 314160 66580 314166 66592
rect 360289 66589 360301 66592
rect 360335 66620 360347 66623
rect 376662 66620 376668 66632
rect 360335 66592 376668 66620
rect 360335 66589 360347 66592
rect 360289 66583 360347 66589
rect 376662 66580 376668 66592
rect 376720 66580 376726 66632
rect 360102 66484 360108 66496
rect 360015 66456 360108 66484
rect 360102 66444 360108 66456
rect 360160 66484 360166 66496
rect 445754 66484 445760 66496
rect 360160 66456 445760 66484
rect 360160 66444 360166 66456
rect 445754 66444 445760 66456
rect 445812 66444 445818 66496
rect 9214 66104 9220 66156
rect 9272 66144 9278 66156
rect 9309 66147 9367 66153
rect 9309 66144 9321 66147
rect 9272 66116 9321 66144
rect 9272 66104 9278 66116
rect 9309 66113 9321 66116
rect 9355 66113 9367 66147
rect 9309 66107 9367 66113
rect 9030 65968 9036 66020
rect 9088 66008 9094 66020
rect 9493 66011 9551 66017
rect 9493 66008 9505 66011
rect 9088 65980 9505 66008
rect 9088 65968 9094 65980
rect 9493 65977 9505 65980
rect 9539 65977 9551 66011
rect 9493 65971 9551 65977
rect 493870 65532 493876 65544
rect 493831 65504 493876 65532
rect 493870 65492 493876 65504
rect 493928 65492 493934 65544
rect 314010 63724 314016 63776
rect 314068 63764 314074 63776
rect 477313 63767 477371 63773
rect 477313 63764 477325 63767
rect 314068 63736 477325 63764
rect 314068 63724 314074 63736
rect 477313 63733 477325 63736
rect 477359 63733 477371 63767
rect 477313 63727 477371 63733
rect 480622 63452 480628 63504
rect 480680 63492 480686 63504
rect 495526 63492 495532 63504
rect 480680 63464 495532 63492
rect 480680 63452 480686 63464
rect 495526 63452 495532 63464
rect 495584 63452 495590 63504
rect 344922 61208 344928 61260
rect 344980 61248 344986 61260
rect 445941 61251 445999 61257
rect 445941 61248 445953 61251
rect 344980 61220 445953 61248
rect 344980 61208 344986 61220
rect 445941 61217 445953 61220
rect 445987 61217 445999 61251
rect 445941 61211 445999 61217
rect 446030 61208 446036 61260
rect 446088 61248 446094 61260
rect 446088 61220 446133 61248
rect 446088 61208 446094 61220
rect 445662 61180 445668 61192
rect 445575 61152 445668 61180
rect 445662 61140 445668 61152
rect 445720 61140 445726 61192
rect 445754 61140 445760 61192
rect 445812 61180 445818 61192
rect 445812 61152 445857 61180
rect 445812 61140 445818 61152
rect 445680 61112 445708 61140
rect 496078 61112 496084 61124
rect 445680 61084 496084 61112
rect 496078 61072 496084 61084
rect 496136 61072 496142 61124
rect 422938 61004 422944 61056
rect 422996 61044 423002 61056
rect 445481 61047 445539 61053
rect 445481 61044 445493 61047
rect 422996 61016 445493 61044
rect 422996 61004 423002 61016
rect 445481 61013 445493 61016
rect 445527 61013 445539 61047
rect 445481 61007 445539 61013
rect 406286 59712 406292 59764
rect 406344 59752 406350 59764
rect 443178 59752 443184 59764
rect 406344 59724 443184 59752
rect 406344 59712 406350 59724
rect 443178 59712 443184 59724
rect 443236 59712 443242 59764
rect 419534 59684 419540 59696
rect 372540 59656 419540 59684
rect 315390 59576 315396 59628
rect 315448 59616 315454 59628
rect 372540 59625 372568 59656
rect 419534 59644 419540 59656
rect 419592 59644 419598 59696
rect 372525 59619 372583 59625
rect 315448 59588 354674 59616
rect 315448 59576 315454 59588
rect 354646 59548 354674 59588
rect 372525 59585 372537 59619
rect 372571 59585 372583 59619
rect 372706 59616 372712 59628
rect 372667 59588 372712 59616
rect 372525 59579 372583 59585
rect 372706 59576 372712 59588
rect 372764 59576 372770 59628
rect 406105 59619 406163 59625
rect 406105 59616 406117 59619
rect 373966 59588 406117 59616
rect 373966 59548 373994 59588
rect 406105 59585 406117 59588
rect 406151 59585 406163 59619
rect 406286 59616 406292 59628
rect 406247 59588 406292 59616
rect 406105 59579 406163 59585
rect 406286 59576 406292 59588
rect 406344 59576 406350 59628
rect 406381 59619 406439 59625
rect 406381 59585 406393 59619
rect 406427 59585 406439 59619
rect 406381 59579 406439 59585
rect 354646 59520 373994 59548
rect 401226 59508 401232 59560
rect 401284 59548 401290 59560
rect 406396 59548 406424 59579
rect 406470 59576 406476 59628
rect 406528 59616 406534 59628
rect 464246 59616 464252 59628
rect 406528 59588 406573 59616
rect 412606 59588 464252 59616
rect 406528 59576 406534 59588
rect 412606 59548 412634 59588
rect 464246 59576 464252 59588
rect 464304 59576 464310 59628
rect 401284 59520 412634 59548
rect 401284 59508 401290 59520
rect 344278 59440 344284 59492
rect 344336 59480 344342 59492
rect 406749 59483 406807 59489
rect 406749 59480 406761 59483
rect 344336 59452 406761 59480
rect 344336 59440 344342 59452
rect 406749 59449 406761 59452
rect 406795 59449 406807 59483
rect 406749 59443 406807 59449
rect 342898 59372 342904 59424
rect 342956 59412 342962 59424
rect 372341 59415 372399 59421
rect 372341 59412 372353 59415
rect 342956 59384 372353 59412
rect 342956 59372 342962 59384
rect 372341 59381 372353 59384
rect 372387 59381 372399 59415
rect 372341 59375 372399 59381
rect 398098 59168 398104 59220
rect 398156 59208 398162 59220
rect 495526 59208 495532 59220
rect 398156 59180 495532 59208
rect 398156 59168 398162 59180
rect 495526 59168 495532 59180
rect 495584 59168 495590 59220
rect 7098 58488 7104 58540
rect 7156 58528 7162 58540
rect 7837 58531 7895 58537
rect 7837 58528 7849 58531
rect 7156 58500 7849 58528
rect 7156 58488 7162 58500
rect 7837 58497 7849 58500
rect 7883 58497 7895 58531
rect 7837 58491 7895 58497
rect 2774 58216 2780 58268
rect 2832 58256 2838 58268
rect 5166 58256 5172 58268
rect 2832 58228 5172 58256
rect 2832 58216 2838 58228
rect 5166 58216 5172 58228
rect 5224 58216 5230 58268
rect 313734 57400 313740 57452
rect 313792 57440 313798 57452
rect 421929 57443 421987 57449
rect 421929 57440 421941 57443
rect 313792 57412 421941 57440
rect 313792 57400 313798 57412
rect 421929 57409 421941 57412
rect 421975 57409 421987 57443
rect 421929 57403 421987 57409
rect 318150 57196 318156 57248
rect 318208 57236 318214 57248
rect 422018 57236 422024 57248
rect 318208 57208 422024 57236
rect 318208 57196 318214 57208
rect 422018 57196 422024 57208
rect 422076 57196 422082 57248
rect 312446 55836 312452 55888
rect 312504 55876 312510 55888
rect 320174 55876 320180 55888
rect 312504 55848 320180 55876
rect 312504 55836 312510 55848
rect 320174 55836 320180 55848
rect 320232 55836 320238 55888
rect 9398 54816 9404 54868
rect 9456 54856 9462 54868
rect 9493 54859 9551 54865
rect 9493 54856 9505 54859
rect 9456 54828 9505 54856
rect 9456 54816 9462 54828
rect 9493 54825 9505 54828
rect 9539 54825 9551 54859
rect 9493 54819 9551 54825
rect 401226 54652 401232 54664
rect 401187 54624 401232 54652
rect 401226 54612 401232 54624
rect 401284 54612 401290 54664
rect 401134 54516 401140 54528
rect 401047 54488 401140 54516
rect 401134 54476 401140 54488
rect 401192 54516 401198 54528
rect 442902 54516 442908 54528
rect 401192 54488 442908 54516
rect 401192 54476 401198 54488
rect 442902 54476 442908 54488
rect 442960 54476 442966 54528
rect 2774 53660 2780 53712
rect 2832 53700 2838 53712
rect 5074 53700 5080 53712
rect 2832 53672 5080 53700
rect 2832 53660 2838 53672
rect 5074 53660 5080 53672
rect 5132 53660 5138 53712
rect 310057 50303 310115 50309
rect 310057 50269 310069 50303
rect 310103 50300 310115 50303
rect 367002 50300 367008 50312
rect 310103 50272 367008 50300
rect 310103 50269 310115 50272
rect 310057 50263 310115 50269
rect 367002 50260 367008 50272
rect 367060 50260 367066 50312
rect 310149 50167 310207 50173
rect 310149 50133 310161 50167
rect 310195 50164 310207 50167
rect 385218 50164 385224 50176
rect 310195 50136 385224 50164
rect 310195 50133 310207 50136
rect 310149 50127 310207 50133
rect 385218 50124 385224 50136
rect 385276 50124 385282 50176
rect 310057 48263 310115 48269
rect 310057 48229 310069 48263
rect 310103 48260 310115 48263
rect 311710 48260 311716 48272
rect 310103 48232 311716 48260
rect 310103 48229 310115 48232
rect 310057 48223 310115 48229
rect 311710 48220 311716 48232
rect 311768 48220 311774 48272
rect 463878 48124 463884 48136
rect 463839 48096 463884 48124
rect 463878 48084 463884 48096
rect 463936 48084 463942 48136
rect 314470 46316 314476 46368
rect 314528 46356 314534 46368
rect 346121 46359 346179 46365
rect 346121 46356 346133 46359
rect 314528 46328 346133 46356
rect 314528 46316 314534 46328
rect 346121 46325 346133 46328
rect 346167 46325 346179 46359
rect 346121 46319 346179 46325
rect 318518 46044 318524 46096
rect 318576 46084 318582 46096
rect 340601 46087 340659 46093
rect 340601 46084 340613 46087
rect 318576 46056 340613 46084
rect 318576 46044 318582 46056
rect 340601 46053 340613 46056
rect 340647 46053 340659 46087
rect 340601 46047 340659 46053
rect 318702 45976 318708 46028
rect 318760 46016 318766 46028
rect 340141 46019 340199 46025
rect 340141 46016 340153 46019
rect 318760 45988 340153 46016
rect 318760 45976 318766 45988
rect 340141 45985 340153 45988
rect 340187 45985 340199 46019
rect 340141 45979 340199 45985
rect 340233 46019 340291 46025
rect 340233 45985 340245 46019
rect 340279 46016 340291 46019
rect 430574 46016 430580 46028
rect 340279 45988 430580 46016
rect 340279 45985 340291 45988
rect 340233 45979 340291 45985
rect 430574 45976 430580 45988
rect 430632 45976 430638 46028
rect 339954 45948 339960 45960
rect 339915 45920 339960 45948
rect 339954 45908 339960 45920
rect 340012 45908 340018 45960
rect 340326 45951 340384 45957
rect 340326 45948 340338 45951
rect 340248 45920 340338 45948
rect 318058 45772 318064 45824
rect 318116 45812 318122 45824
rect 339865 45815 339923 45821
rect 339865 45812 339877 45815
rect 318116 45784 339877 45812
rect 318116 45772 318122 45784
rect 339865 45781 339877 45784
rect 339911 45781 339923 45815
rect 340248 45812 340276 45920
rect 340326 45917 340338 45920
rect 340372 45917 340384 45951
rect 340326 45911 340384 45917
rect 340509 45951 340567 45957
rect 340509 45917 340521 45951
rect 340555 45948 340567 45951
rect 340601 45951 340659 45957
rect 340601 45948 340613 45951
rect 340555 45920 340613 45948
rect 340555 45917 340567 45920
rect 340509 45911 340567 45917
rect 340601 45917 340613 45920
rect 340647 45917 340659 45951
rect 498197 45951 498255 45957
rect 498197 45948 498209 45951
rect 340601 45911 340659 45917
rect 344986 45920 498209 45948
rect 340414 45812 340420 45824
rect 340248 45784 340420 45812
rect 339865 45775 339923 45781
rect 340414 45772 340420 45784
rect 340472 45812 340478 45824
rect 344986 45812 345014 45920
rect 498197 45917 498209 45920
rect 498243 45917 498255 45951
rect 498197 45911 498255 45917
rect 340472 45784 345014 45812
rect 340472 45772 340478 45784
rect 369210 45500 369216 45552
rect 369268 45540 369274 45552
rect 495526 45540 495532 45552
rect 369268 45512 495532 45540
rect 369268 45500 369274 45512
rect 495526 45500 495532 45512
rect 495584 45500 495590 45552
rect 310057 45067 310115 45073
rect 310057 45033 310069 45067
rect 310103 45064 310115 45067
rect 311894 45064 311900 45076
rect 310103 45036 311900 45064
rect 310103 45033 310115 45036
rect 310057 45027 310115 45033
rect 311894 45024 311900 45036
rect 311952 45024 311958 45076
rect 310146 44888 310152 44940
rect 310204 44928 310210 44940
rect 310609 44931 310667 44937
rect 310609 44928 310621 44931
rect 310204 44900 310621 44928
rect 310204 44888 310210 44900
rect 310609 44897 310621 44900
rect 310655 44928 310667 44931
rect 378962 44928 378968 44940
rect 310655 44900 378968 44928
rect 310655 44897 310667 44900
rect 310609 44891 310667 44897
rect 378962 44888 378968 44900
rect 379020 44888 379026 44940
rect 310422 44860 310428 44872
rect 310383 44832 310428 44860
rect 310422 44820 310428 44832
rect 310480 44820 310486 44872
rect 310238 44684 310244 44736
rect 310296 44724 310302 44736
rect 310517 44727 310575 44733
rect 310517 44724 310529 44727
rect 310296 44696 310529 44724
rect 310296 44684 310302 44696
rect 310517 44693 310529 44696
rect 310563 44693 310575 44727
rect 310517 44687 310575 44693
rect 310241 43095 310299 43101
rect 310241 43061 310253 43095
rect 310287 43092 310299 43095
rect 496354 43092 496360 43104
rect 310287 43064 496360 43092
rect 310287 43061 310299 43064
rect 310241 43055 310299 43061
rect 496354 43052 496360 43064
rect 496412 43052 496418 43104
rect 8288 42279 8346 42285
rect 8288 42245 8300 42279
rect 8334 42276 8346 42279
rect 8386 42276 8392 42288
rect 8334 42248 8392 42276
rect 8334 42245 8346 42248
rect 8288 42239 8346 42245
rect 8386 42236 8392 42248
rect 8444 42236 8450 42288
rect 8018 42140 8024 42152
rect 7979 42112 8024 42140
rect 8018 42100 8024 42112
rect 8076 42100 8082 42152
rect 9398 42004 9404 42016
rect 9359 41976 9404 42004
rect 9398 41964 9404 41976
rect 9456 41964 9462 42016
rect 338758 39788 338764 39840
rect 338816 39828 338822 39840
rect 366821 39831 366879 39837
rect 366821 39828 366833 39831
rect 338816 39800 366833 39828
rect 338816 39788 338822 39800
rect 366821 39797 366833 39800
rect 366867 39797 366879 39831
rect 366821 39791 366879 39797
rect 384298 37816 384304 37868
rect 384356 37856 384362 37868
rect 418249 37859 418307 37865
rect 418249 37856 418261 37859
rect 384356 37828 418261 37856
rect 384356 37816 384362 37828
rect 418249 37825 418261 37828
rect 418295 37825 418307 37859
rect 418249 37819 418307 37825
rect 418338 37788 418344 37800
rect 418299 37760 418344 37788
rect 418338 37748 418344 37760
rect 418396 37748 418402 37800
rect 418430 37748 418436 37800
rect 418488 37788 418494 37800
rect 479426 37788 479432 37800
rect 418488 37760 479432 37788
rect 418488 37748 418494 37760
rect 479426 37748 479432 37760
rect 479484 37748 479490 37800
rect 310241 37655 310299 37661
rect 310241 37621 310253 37655
rect 310287 37652 310299 37655
rect 395338 37652 395344 37664
rect 310287 37624 395344 37652
rect 310287 37621 310299 37624
rect 310241 37615 310299 37621
rect 395338 37612 395344 37624
rect 395396 37612 395402 37664
rect 417878 37652 417884 37664
rect 417839 37624 417884 37652
rect 417878 37612 417884 37624
rect 417936 37612 417942 37664
rect 312722 36660 312728 36712
rect 312780 36700 312786 36712
rect 368474 36700 368480 36712
rect 312780 36672 368480 36700
rect 312780 36660 312786 36672
rect 368474 36660 368480 36672
rect 368532 36660 368538 36712
rect 312630 36592 312636 36644
rect 312688 36632 312694 36644
rect 463878 36632 463884 36644
rect 312688 36604 463884 36632
rect 312688 36592 312694 36604
rect 463878 36592 463884 36604
rect 463936 36592 463942 36644
rect 311618 36524 311624 36576
rect 311676 36564 311682 36576
rect 466454 36564 466460 36576
rect 311676 36536 466460 36564
rect 311676 36524 311682 36536
rect 466454 36524 466460 36536
rect 466512 36524 466518 36576
rect 342533 36363 342591 36369
rect 342533 36329 342545 36363
rect 342579 36360 342591 36363
rect 346486 36360 346492 36372
rect 342579 36332 346492 36360
rect 342579 36329 342591 36332
rect 342533 36323 342591 36329
rect 346486 36320 346492 36332
rect 346544 36320 346550 36372
rect 343910 36156 343916 36168
rect 343871 36128 343916 36156
rect 343910 36116 343916 36128
rect 343968 36156 343974 36168
rect 373166 36156 373172 36168
rect 343968 36128 373172 36156
rect 343968 36116 343974 36128
rect 373166 36116 373172 36128
rect 373224 36116 373230 36168
rect 343668 36091 343726 36097
rect 343668 36057 343680 36091
rect 343714 36088 343726 36091
rect 346302 36088 346308 36100
rect 343714 36060 346308 36088
rect 343714 36057 343726 36060
rect 343668 36051 343726 36057
rect 346302 36048 346308 36060
rect 346360 36048 346366 36100
rect 410518 35844 410524 35896
rect 410576 35884 410582 35896
rect 495526 35884 495532 35896
rect 410576 35856 495532 35884
rect 410576 35844 410582 35856
rect 495526 35844 495532 35856
rect 495584 35844 495590 35896
rect 390922 35272 390928 35284
rect 390883 35244 390928 35272
rect 390922 35232 390928 35244
rect 390980 35232 390986 35284
rect 392026 35068 392032 35080
rect 392084 35077 392090 35080
rect 391996 35040 392032 35068
rect 392026 35028 392032 35040
rect 392084 35031 392096 35077
rect 392305 35071 392363 35077
rect 392305 35037 392317 35071
rect 392351 35068 392363 35071
rect 392489 35071 392547 35077
rect 392489 35068 392501 35071
rect 392351 35040 392501 35068
rect 392351 35037 392363 35040
rect 392305 35031 392363 35037
rect 392489 35037 392501 35040
rect 392535 35068 392547 35071
rect 416866 35068 416872 35080
rect 392535 35040 416872 35068
rect 392535 35037 392547 35040
rect 392489 35031 392547 35037
rect 392084 35028 392090 35031
rect 416866 35028 416872 35040
rect 416924 35028 416930 35080
rect 371786 34728 371792 34740
rect 371747 34700 371792 34728
rect 371786 34688 371792 34700
rect 371844 34688 371850 34740
rect 372890 34592 372896 34604
rect 372948 34601 372954 34604
rect 372860 34564 372896 34592
rect 372890 34552 372896 34564
rect 372948 34555 372960 34601
rect 373166 34592 373172 34604
rect 373127 34564 373172 34592
rect 372948 34552 372954 34555
rect 373166 34552 373172 34564
rect 373224 34592 373230 34604
rect 373224 34564 373994 34592
rect 373224 34552 373230 34564
rect 373966 34524 373994 34564
rect 392489 34527 392547 34533
rect 392489 34524 392501 34527
rect 373966 34496 392501 34524
rect 392489 34493 392501 34496
rect 392535 34493 392547 34527
rect 392489 34487 392547 34493
rect 399478 32008 399484 32020
rect 399439 31980 399484 32008
rect 399478 31968 399484 31980
rect 399536 31968 399542 32020
rect 321370 31424 321376 31476
rect 321428 31464 321434 31476
rect 416682 31464 416688 31476
rect 321428 31436 412634 31464
rect 321428 31424 321434 31436
rect 412606 31328 412634 31436
rect 416608 31436 416688 31464
rect 416608 31405 416636 31436
rect 416682 31424 416688 31436
rect 416740 31424 416746 31476
rect 417510 31464 417516 31476
rect 417471 31436 417516 31464
rect 417510 31424 417516 31436
rect 417568 31424 417574 31476
rect 416602 31399 416660 31405
rect 416602 31365 416614 31399
rect 416648 31365 416660 31399
rect 416602 31359 416660 31365
rect 416866 31356 416872 31408
rect 416924 31396 416930 31408
rect 416924 31368 418936 31396
rect 416924 31356 416930 31368
rect 418908 31337 418936 31368
rect 418626 31331 418684 31337
rect 418626 31328 418638 31331
rect 412606 31300 418638 31328
rect 418626 31297 418638 31300
rect 418672 31297 418684 31331
rect 418626 31291 418684 31297
rect 418893 31331 418951 31337
rect 418893 31297 418905 31331
rect 418939 31328 418951 31331
rect 418939 31300 422294 31328
rect 418939 31297 418951 31300
rect 418893 31291 418951 31297
rect 416866 31260 416872 31272
rect 416827 31232 416872 31260
rect 416866 31220 416872 31232
rect 416924 31220 416930 31272
rect 422266 31260 422294 31300
rect 458174 31260 458180 31272
rect 422266 31232 458180 31260
rect 458174 31220 458180 31232
rect 458232 31220 458238 31272
rect 415486 31124 415492 31136
rect 415399 31096 415492 31124
rect 415486 31084 415492 31096
rect 415544 31124 415550 31136
rect 463510 31124 463516 31136
rect 415544 31096 463516 31124
rect 415544 31084 415550 31096
rect 463510 31084 463516 31096
rect 463568 31084 463574 31136
rect 311342 30676 311348 30728
rect 311400 30716 311406 30728
rect 408497 30719 408555 30725
rect 408497 30716 408509 30719
rect 311400 30688 408509 30716
rect 311400 30676 311406 30688
rect 408497 30685 408509 30688
rect 408543 30685 408555 30719
rect 408497 30679 408555 30685
rect 318334 30268 318340 30320
rect 318392 30308 318398 30320
rect 320450 30308 320456 30320
rect 318392 30280 320456 30308
rect 318392 30268 318398 30280
rect 320450 30268 320456 30280
rect 320508 30268 320514 30320
rect 318426 30200 318432 30252
rect 318484 30240 318490 30252
rect 320361 30243 320419 30249
rect 320361 30240 320373 30243
rect 318484 30212 320373 30240
rect 318484 30200 318490 30212
rect 320361 30209 320373 30212
rect 320407 30209 320419 30243
rect 320361 30203 320419 30209
rect 376018 27452 376024 27464
rect 375979 27424 376024 27452
rect 376018 27412 376024 27424
rect 376076 27412 376082 27464
rect 9306 25888 9312 25900
rect 9267 25860 9312 25888
rect 9306 25848 9312 25860
rect 9364 25848 9370 25900
rect 9490 25820 9496 25832
rect 9451 25792 9496 25820
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 9125 25687 9183 25693
rect 9125 25653 9137 25687
rect 9171 25684 9183 25687
rect 9214 25684 9220 25696
rect 9171 25656 9220 25684
rect 9171 25653 9183 25656
rect 9125 25647 9183 25653
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 310146 25344 310152 25356
rect 310107 25316 310152 25344
rect 310146 25304 310152 25316
rect 310204 25304 310210 25356
rect 310333 25347 310391 25353
rect 310333 25313 310345 25347
rect 310379 25344 310391 25347
rect 310606 25344 310612 25356
rect 310379 25316 310612 25344
rect 310379 25313 310391 25316
rect 310333 25307 310391 25313
rect 310606 25304 310612 25316
rect 310664 25304 310670 25356
rect 310425 25279 310483 25285
rect 310425 25245 310437 25279
rect 310471 25276 310483 25279
rect 311526 25276 311532 25288
rect 310471 25248 311532 25276
rect 310471 25245 310483 25248
rect 310425 25239 310483 25245
rect 311526 25236 311532 25248
rect 311584 25236 311590 25288
rect 310793 25143 310851 25149
rect 310793 25109 310805 25143
rect 310839 25140 310851 25143
rect 360194 25140 360200 25152
rect 310839 25112 360200 25140
rect 310839 25109 310851 25112
rect 310793 25103 310851 25109
rect 360194 25100 360200 25112
rect 360252 25100 360258 25152
rect 356698 23400 356704 23452
rect 356756 23440 356762 23452
rect 495526 23440 495532 23452
rect 356756 23412 495532 23440
rect 356756 23400 356762 23412
rect 495526 23400 495532 23412
rect 495584 23400 495590 23452
rect 456058 16096 456064 16108
rect 456019 16068 456064 16096
rect 456058 16056 456064 16068
rect 456116 16056 456122 16108
rect 317138 15852 317144 15904
rect 317196 15892 317202 15904
rect 455877 15895 455935 15901
rect 455877 15892 455889 15895
rect 317196 15864 455889 15892
rect 317196 15852 317202 15864
rect 455877 15861 455889 15864
rect 455923 15861 455935 15895
rect 455877 15855 455935 15861
rect 318242 15444 318248 15496
rect 318300 15484 318306 15496
rect 335415 15487 335473 15493
rect 335415 15484 335427 15487
rect 318300 15456 335427 15484
rect 318300 15444 318306 15456
rect 335415 15453 335427 15456
rect 335461 15453 335473 15487
rect 335633 15487 335691 15493
rect 335415 15447 335473 15453
rect 335540 15465 335598 15471
rect 335540 15431 335552 15465
rect 335586 15431 335598 15465
rect 335633 15453 335645 15487
rect 335679 15453 335691 15487
rect 335633 15447 335691 15453
rect 335817 15487 335875 15493
rect 335817 15453 335829 15487
rect 335863 15484 335875 15487
rect 453022 15484 453028 15496
rect 335863 15456 453028 15484
rect 335863 15453 335875 15456
rect 335817 15447 335875 15453
rect 315666 15376 315672 15428
rect 315724 15416 315730 15428
rect 335540 15425 335598 15431
rect 335173 15419 335231 15425
rect 335173 15416 335185 15419
rect 315724 15388 335185 15416
rect 315724 15376 315730 15388
rect 335173 15385 335185 15388
rect 335219 15385 335231 15419
rect 335173 15379 335231 15385
rect 335556 15360 335584 15425
rect 335648 15360 335676 15447
rect 453022 15444 453028 15456
rect 453080 15444 453086 15496
rect 496354 15484 496360 15496
rect 496315 15456 496360 15484
rect 496354 15444 496360 15456
rect 496412 15444 496418 15496
rect 335538 15308 335544 15360
rect 335596 15308 335602 15360
rect 335630 15308 335636 15360
rect 335688 15308 335694 15360
rect 447778 15308 447784 15360
rect 447836 15348 447842 15360
rect 496449 15351 496507 15357
rect 496449 15348 496461 15351
rect 447836 15320 496461 15348
rect 447836 15308 447842 15320
rect 496449 15317 496461 15320
rect 496495 15317 496507 15351
rect 496449 15311 496507 15317
rect 475378 14016 475384 14068
rect 475436 14056 475442 14068
rect 479245 14059 479303 14065
rect 479245 14056 479257 14059
rect 475436 14028 479257 14056
rect 475436 14016 475442 14028
rect 479245 14025 479257 14028
rect 479291 14025 479303 14059
rect 479245 14019 479303 14025
rect 460198 13948 460204 14000
rect 460256 13988 460262 14000
rect 479337 13991 479395 13997
rect 479337 13988 479349 13991
rect 460256 13960 479349 13988
rect 460256 13948 460262 13960
rect 479337 13957 479349 13960
rect 479383 13957 479395 13991
rect 479337 13951 479395 13957
rect 414658 13812 414664 13864
rect 414716 13852 414722 13864
rect 478785 13855 478843 13861
rect 478785 13852 478797 13855
rect 414716 13824 478797 13852
rect 414716 13812 414722 13824
rect 478785 13821 478797 13824
rect 478831 13821 478843 13855
rect 478785 13815 478843 13821
rect 479426 13812 479432 13864
rect 479484 13852 479490 13864
rect 479484 13824 479529 13852
rect 479484 13812 479490 13824
rect 351178 13744 351184 13796
rect 351236 13784 351242 13796
rect 495434 13784 495440 13796
rect 351236 13756 495440 13784
rect 351236 13744 351242 13756
rect 495434 13744 495440 13756
rect 495492 13744 495498 13796
rect 478785 13719 478843 13725
rect 478785 13685 478797 13719
rect 478831 13716 478843 13719
rect 478877 13719 478935 13725
rect 478877 13716 478889 13719
rect 478831 13688 478889 13716
rect 478831 13685 478843 13688
rect 478785 13679 478843 13685
rect 478877 13685 478889 13688
rect 478923 13685 478935 13719
rect 478877 13679 478935 13685
rect 344646 12424 344652 12436
rect 344607 12396 344652 12424
rect 344646 12384 344652 12396
rect 344704 12384 344710 12436
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 417878 11880 417884 11892
rect 9548 11852 417884 11880
rect 9548 11840 9554 11852
rect 417878 11840 417884 11852
rect 417936 11840 417942 11892
rect 261846 10616 261852 10668
rect 261904 10656 261910 10668
rect 315482 10656 315488 10668
rect 261904 10628 315488 10656
rect 261904 10616 261910 10628
rect 315482 10616 315488 10628
rect 315540 10616 315546 10668
rect 239950 10548 239956 10600
rect 240008 10588 240014 10600
rect 310146 10588 310152 10600
rect 240008 10560 310152 10588
rect 240008 10548 240014 10560
rect 310146 10548 310152 10560
rect 310204 10548 310210 10600
rect 244642 10480 244648 10532
rect 244700 10520 244706 10532
rect 450262 10520 450268 10532
rect 244700 10492 450268 10520
rect 244700 10480 244706 10492
rect 450262 10480 450268 10492
rect 450320 10480 450326 10532
rect 147950 10412 147956 10464
rect 148008 10452 148014 10464
rect 371786 10452 371792 10464
rect 148008 10424 371792 10452
rect 148008 10412 148014 10424
rect 371786 10412 371792 10424
rect 371844 10412 371850 10464
rect 116762 10344 116768 10396
rect 116820 10384 116826 10396
rect 342346 10384 342352 10396
rect 116820 10356 342352 10384
rect 116820 10344 116826 10356
rect 342346 10344 342352 10356
rect 342404 10344 342410 10396
rect 151262 10276 151268 10328
rect 151320 10316 151326 10328
rect 383746 10316 383752 10328
rect 151320 10288 383752 10316
rect 151320 10276 151326 10288
rect 383746 10276 383752 10288
rect 383804 10276 383810 10328
rect 168650 9868 168656 9920
rect 168708 9908 168714 9920
rect 169110 9908 169116 9920
rect 168708 9880 169116 9908
rect 168708 9868 168714 9880
rect 169110 9868 169116 9880
rect 169168 9868 169174 9920
rect 278133 9911 278191 9917
rect 278133 9908 278145 9911
rect 277596 9880 278145 9908
rect 78217 9707 78275 9713
rect 78217 9673 78229 9707
rect 78263 9673 78275 9707
rect 151262 9704 151268 9716
rect 151223 9676 151268 9704
rect 78217 9667 78275 9673
rect 77294 9596 77300 9648
rect 77352 9636 77358 9648
rect 78232 9636 78260 9667
rect 151262 9664 151268 9676
rect 151320 9664 151326 9716
rect 168650 9664 168656 9716
rect 168708 9704 168714 9716
rect 168708 9676 168788 9704
rect 168708 9664 168714 9676
rect 78582 9636 78588 9648
rect 77352 9608 78076 9636
rect 78232 9608 78588 9636
rect 77352 9596 77358 9608
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 35345 9571 35403 9577
rect 35345 9568 35357 9571
rect 8812 9540 35357 9568
rect 8812 9528 8818 9540
rect 35345 9537 35357 9540
rect 35391 9568 35403 9571
rect 35713 9571 35771 9577
rect 35713 9568 35725 9571
rect 35391 9540 35725 9568
rect 35391 9537 35403 9540
rect 35345 9531 35403 9537
rect 35713 9537 35725 9540
rect 35759 9537 35771 9571
rect 35713 9531 35771 9537
rect 65337 9571 65395 9577
rect 65337 9537 65349 9571
rect 65383 9568 65395 9571
rect 66165 9571 66223 9577
rect 66165 9568 66177 9571
rect 65383 9540 66177 9568
rect 65383 9537 65395 9540
rect 65337 9531 65395 9537
rect 66165 9537 66177 9540
rect 66211 9537 66223 9571
rect 77110 9568 77116 9580
rect 77071 9540 77116 9568
rect 66165 9531 66223 9537
rect 77110 9528 77116 9540
rect 77168 9528 77174 9580
rect 77205 9571 77263 9577
rect 77205 9537 77217 9571
rect 77251 9568 77263 9571
rect 77481 9571 77539 9577
rect 77481 9568 77493 9571
rect 77251 9540 77493 9568
rect 77251 9537 77263 9540
rect 77205 9531 77263 9537
rect 77481 9537 77493 9540
rect 77527 9537 77539 9571
rect 77846 9568 77852 9580
rect 77807 9540 77852 9568
rect 77481 9531 77539 9537
rect 77846 9528 77852 9540
rect 77904 9528 77910 9580
rect 78048 9577 78076 9608
rect 78582 9596 78588 9608
rect 78640 9596 78646 9648
rect 168760 9636 168788 9676
rect 168926 9674 168932 9716
rect 168852 9664 168932 9674
rect 168984 9664 168990 9716
rect 185397 9707 185455 9713
rect 169110 9674 169116 9686
rect 168852 9648 168972 9664
rect 78784 9608 168788 9636
rect 78033 9571 78091 9577
rect 78033 9537 78045 9571
rect 78079 9537 78091 9571
rect 78033 9531 78091 9537
rect 78401 9571 78459 9577
rect 78401 9537 78413 9571
rect 78447 9568 78459 9571
rect 78784 9568 78812 9608
rect 168834 9596 168840 9648
rect 168892 9646 168972 9648
rect 169061 9646 169116 9674
rect 168892 9596 168898 9646
rect 169110 9634 169116 9646
rect 169168 9636 169174 9686
rect 185397 9673 185409 9707
rect 185443 9704 185455 9707
rect 186225 9707 186283 9713
rect 186225 9704 186237 9707
rect 185443 9676 186237 9704
rect 185443 9673 185455 9676
rect 185397 9667 185455 9673
rect 186225 9673 186237 9676
rect 186271 9673 186283 9707
rect 239950 9704 239956 9716
rect 239911 9676 239956 9704
rect 186225 9667 186283 9673
rect 239950 9664 239956 9676
rect 240008 9664 240014 9716
rect 248138 9704 248144 9716
rect 248099 9676 248144 9704
rect 248138 9664 248144 9676
rect 248196 9664 248202 9716
rect 270957 9707 271015 9713
rect 270957 9673 270969 9707
rect 271003 9704 271015 9707
rect 271509 9707 271567 9713
rect 271509 9704 271521 9707
rect 271003 9676 271521 9704
rect 271003 9673 271015 9676
rect 270957 9667 271015 9673
rect 271509 9673 271521 9676
rect 271555 9673 271567 9707
rect 271509 9667 271567 9673
rect 272334 9664 272340 9716
rect 272392 9674 272398 9716
rect 277596 9704 277624 9880
rect 278133 9877 278145 9880
rect 278179 9877 278191 9911
rect 278133 9871 278191 9877
rect 277762 9704 277768 9716
rect 277504 9676 277624 9704
rect 277675 9676 277768 9704
rect 272392 9664 272472 9674
rect 272150 9636 272156 9648
rect 169168 9634 272156 9636
rect 169128 9608 272156 9634
rect 272150 9596 272156 9608
rect 272208 9596 272214 9648
rect 272352 9646 272472 9664
rect 78447 9540 78812 9568
rect 78447 9537 78459 9540
rect 78401 9531 78459 9537
rect 78858 9528 78864 9580
rect 78916 9568 78922 9580
rect 78916 9540 78961 9568
rect 78916 9528 78922 9540
rect 79042 9528 79048 9580
rect 79100 9568 79106 9580
rect 88426 9568 88432 9580
rect 79100 9540 79145 9568
rect 88387 9540 88432 9568
rect 79100 9528 79106 9540
rect 88426 9528 88432 9540
rect 88484 9528 88490 9580
rect 88610 9568 88616 9580
rect 88571 9540 88616 9568
rect 88610 9528 88616 9540
rect 88668 9528 88674 9580
rect 95142 9568 95148 9580
rect 95103 9540 95148 9568
rect 95142 9528 95148 9540
rect 95200 9528 95206 9580
rect 115845 9571 115903 9577
rect 115845 9537 115857 9571
rect 115891 9568 115903 9571
rect 116486 9568 116492 9580
rect 115891 9540 116348 9568
rect 116447 9540 116492 9568
rect 115891 9537 115903 9540
rect 115845 9531 115903 9537
rect 79226 9500 79232 9512
rect 64846 9472 79088 9500
rect 79187 9472 79232 9500
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 64846 9432 64874 9472
rect 65150 9432 65156 9444
rect 7800 9404 64874 9432
rect 65111 9404 65156 9432
rect 7800 9392 7806 9404
rect 65150 9392 65156 9404
rect 65208 9392 65214 9444
rect 76745 9435 76803 9441
rect 76745 9401 76757 9435
rect 76791 9432 76803 9435
rect 77021 9435 77079 9441
rect 77021 9432 77033 9435
rect 76791 9404 77033 9432
rect 76791 9401 76803 9404
rect 76745 9395 76803 9401
rect 77021 9401 77033 9404
rect 77067 9401 77079 9435
rect 79060 9432 79088 9472
rect 79226 9460 79232 9472
rect 79284 9460 79290 9512
rect 116029 9503 116087 9509
rect 103486 9472 115980 9500
rect 88334 9432 88340 9444
rect 79060 9404 84194 9432
rect 88295 9404 88340 9432
rect 77021 9395 77079 9401
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 4798 9364 4804 9376
rect 2832 9336 4804 9364
rect 2832 9324 2838 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 35526 9364 35532 9376
rect 35487 9336 35532 9364
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 72234 9364 72240 9376
rect 72195 9336 72240 9364
rect 72234 9324 72240 9336
rect 72292 9324 72298 9376
rect 77938 9364 77944 9376
rect 77899 9336 77944 9364
rect 77938 9324 77944 9336
rect 77996 9324 78002 9376
rect 84166 9364 84194 9404
rect 88334 9392 88340 9404
rect 88392 9392 88398 9444
rect 103486 9432 103514 9472
rect 93826 9404 103514 9432
rect 115952 9432 115980 9472
rect 116029 9469 116041 9503
rect 116075 9500 116087 9503
rect 116213 9503 116271 9509
rect 116213 9500 116225 9503
rect 116075 9472 116225 9500
rect 116075 9469 116087 9472
rect 116029 9463 116087 9469
rect 116213 9469 116225 9472
rect 116259 9469 116271 9503
rect 116320 9500 116348 9540
rect 116486 9528 116492 9540
rect 116544 9528 116550 9580
rect 116578 9528 116584 9580
rect 116636 9568 116642 9580
rect 116762 9568 116768 9580
rect 116636 9540 116681 9568
rect 116723 9540 116768 9568
rect 116636 9528 116642 9540
rect 116762 9528 116768 9540
rect 116820 9528 116826 9580
rect 147950 9568 147956 9580
rect 147911 9540 147956 9568
rect 147950 9528 147956 9540
rect 148008 9528 148014 9580
rect 148042 9528 148048 9580
rect 148100 9568 148106 9580
rect 150986 9568 150992 9580
rect 148100 9540 148145 9568
rect 148244 9540 150848 9568
rect 150947 9540 150992 9568
rect 148100 9528 148106 9540
rect 121457 9503 121515 9509
rect 121457 9500 121469 9503
rect 116320 9472 121469 9500
rect 116213 9463 116271 9469
rect 121457 9469 121469 9472
rect 121503 9469 121515 9503
rect 121457 9463 121515 9469
rect 138017 9503 138075 9509
rect 138017 9469 138029 9503
rect 138063 9500 138075 9503
rect 138385 9503 138443 9509
rect 138385 9500 138397 9503
rect 138063 9472 138397 9500
rect 138063 9469 138075 9472
rect 138017 9463 138075 9469
rect 138385 9469 138397 9472
rect 138431 9469 138443 9503
rect 148244 9500 148272 9540
rect 138385 9463 138443 9469
rect 146864 9472 148272 9500
rect 148321 9503 148379 9509
rect 142157 9435 142215 9441
rect 142157 9432 142169 9435
rect 115952 9404 142169 9432
rect 93826 9364 93854 9404
rect 142157 9401 142169 9404
rect 142203 9401 142215 9435
rect 142157 9395 142215 9401
rect 98822 9364 98828 9376
rect 84166 9336 93854 9364
rect 98783 9336 98828 9364
rect 98822 9324 98828 9336
rect 98880 9324 98886 9376
rect 111705 9367 111763 9373
rect 111705 9333 111717 9367
rect 111751 9364 111763 9367
rect 115845 9367 115903 9373
rect 115845 9364 115857 9367
rect 111751 9336 115857 9364
rect 111751 9333 111763 9336
rect 111705 9327 111763 9333
rect 115845 9333 115857 9336
rect 115891 9333 115903 9367
rect 115845 9327 115903 9333
rect 115937 9367 115995 9373
rect 115937 9333 115949 9367
rect 115983 9364 115995 9367
rect 116305 9367 116363 9373
rect 116305 9364 116317 9367
rect 115983 9336 116317 9364
rect 115983 9333 115995 9336
rect 115937 9327 115995 9333
rect 116305 9333 116317 9336
rect 116351 9333 116363 9367
rect 116305 9327 116363 9333
rect 120077 9367 120135 9373
rect 120077 9333 120089 9367
rect 120123 9364 120135 9367
rect 121181 9367 121239 9373
rect 121181 9364 121193 9367
rect 120123 9336 121193 9364
rect 120123 9333 120135 9336
rect 120077 9327 120135 9333
rect 121181 9333 121193 9336
rect 121227 9333 121239 9367
rect 121181 9327 121239 9333
rect 121457 9367 121515 9373
rect 121457 9333 121469 9367
rect 121503 9364 121515 9367
rect 146864 9364 146892 9472
rect 148321 9469 148333 9503
rect 148367 9500 148379 9503
rect 148965 9503 149023 9509
rect 148965 9500 148977 9503
rect 148367 9472 148977 9500
rect 148367 9469 148379 9472
rect 148321 9463 148379 9469
rect 148965 9469 148977 9472
rect 149011 9469 149023 9503
rect 148965 9463 149023 9469
rect 150529 9503 150587 9509
rect 150529 9469 150541 9503
rect 150575 9500 150587 9503
rect 150713 9503 150771 9509
rect 150713 9500 150725 9503
rect 150575 9472 150725 9500
rect 150575 9469 150587 9472
rect 150529 9463 150587 9469
rect 150713 9469 150725 9472
rect 150759 9469 150771 9503
rect 150820 9500 150848 9540
rect 150986 9528 150992 9540
rect 151044 9528 151050 9580
rect 151081 9571 151139 9577
rect 151081 9537 151093 9571
rect 151127 9568 151139 9571
rect 151725 9571 151783 9577
rect 151725 9568 151737 9571
rect 151127 9540 151737 9568
rect 151127 9537 151139 9540
rect 151081 9531 151139 9537
rect 151725 9537 151737 9540
rect 151771 9537 151783 9571
rect 152550 9568 152556 9580
rect 152511 9540 152556 9568
rect 151725 9531 151783 9537
rect 152550 9528 152556 9540
rect 152608 9528 152614 9580
rect 152737 9571 152795 9577
rect 152737 9537 152749 9571
rect 152783 9568 152795 9571
rect 152921 9571 152979 9577
rect 152921 9568 152933 9571
rect 152783 9540 152933 9568
rect 152783 9537 152795 9540
rect 152737 9531 152795 9537
rect 152921 9537 152933 9540
rect 152967 9537 152979 9571
rect 168742 9568 168748 9580
rect 152921 9531 152979 9537
rect 161446 9540 168748 9568
rect 153013 9503 153071 9509
rect 150820 9472 152596 9500
rect 150713 9463 150771 9469
rect 152461 9435 152519 9441
rect 152461 9432 152473 9435
rect 121503 9336 146892 9364
rect 147048 9404 152473 9432
rect 121503 9333 121515 9336
rect 121457 9327 121515 9333
rect 142157 9299 142215 9305
rect 142157 9265 142169 9299
rect 142203 9296 142215 9299
rect 147048 9296 147076 9404
rect 152461 9401 152473 9404
rect 152507 9401 152519 9435
rect 152568 9432 152596 9472
rect 153013 9469 153025 9503
rect 153059 9500 153071 9503
rect 161446 9500 161474 9540
rect 168742 9528 168748 9540
rect 168800 9528 168806 9580
rect 168926 9577 168932 9580
rect 168920 9568 168932 9577
rect 168887 9540 168932 9568
rect 168920 9531 168932 9540
rect 168926 9528 168932 9531
rect 168984 9528 168990 9580
rect 169294 9528 169300 9580
rect 169352 9568 169358 9580
rect 185489 9571 185547 9577
rect 169352 9540 176654 9568
rect 169352 9528 169358 9540
rect 168650 9500 168656 9512
rect 153059 9472 161474 9500
rect 168611 9472 168656 9500
rect 153059 9469 153071 9472
rect 153013 9463 153071 9469
rect 168650 9460 168656 9472
rect 168708 9460 168714 9512
rect 176626 9500 176654 9540
rect 185489 9537 185501 9571
rect 185535 9568 185547 9571
rect 191193 9571 191251 9577
rect 191193 9568 191205 9571
rect 185535 9540 191205 9568
rect 185535 9537 185547 9540
rect 185489 9531 185547 9537
rect 191193 9537 191205 9540
rect 191239 9537 191251 9571
rect 239858 9568 239864 9580
rect 239819 9540 239864 9568
rect 191193 9531 191251 9537
rect 239858 9528 239864 9540
rect 239916 9528 239922 9580
rect 240042 9568 240048 9580
rect 240003 9540 240048 9568
rect 240042 9528 240048 9540
rect 240100 9528 240106 9580
rect 241517 9571 241575 9577
rect 241517 9537 241529 9571
rect 241563 9568 241575 9571
rect 244550 9568 244556 9580
rect 241563 9540 244412 9568
rect 244511 9540 244556 9568
rect 241563 9537 241575 9540
rect 241517 9531 241575 9537
rect 244274 9500 244280 9512
rect 176626 9472 243584 9500
rect 244235 9472 244280 9500
rect 233881 9435 233939 9441
rect 152568 9404 168696 9432
rect 152461 9395 152519 9401
rect 147766 9364 147772 9376
rect 147727 9336 147772 9364
rect 147766 9324 147772 9336
rect 147824 9324 147830 9376
rect 148229 9367 148287 9373
rect 148229 9333 148241 9367
rect 148275 9364 148287 9367
rect 148505 9367 148563 9373
rect 148505 9364 148517 9367
rect 148275 9336 148517 9364
rect 148275 9333 148287 9336
rect 148229 9327 148287 9333
rect 148505 9333 148517 9336
rect 148551 9333 148563 9367
rect 148505 9327 148563 9333
rect 150437 9367 150495 9373
rect 150437 9333 150449 9367
rect 150483 9364 150495 9367
rect 150805 9367 150863 9373
rect 150805 9364 150817 9367
rect 150483 9336 150817 9364
rect 150483 9333 150495 9336
rect 150437 9327 150495 9333
rect 150805 9333 150817 9336
rect 150851 9333 150863 9367
rect 150805 9327 150863 9333
rect 151725 9367 151783 9373
rect 151725 9333 151737 9367
rect 151771 9364 151783 9367
rect 161477 9367 161535 9373
rect 151771 9336 157334 9364
rect 151771 9333 151783 9336
rect 151725 9327 151783 9333
rect 142203 9268 147076 9296
rect 157306 9296 157334 9336
rect 161477 9333 161489 9367
rect 161523 9364 161535 9367
rect 168377 9367 168435 9373
rect 168377 9364 168389 9367
rect 161523 9336 168389 9364
rect 161523 9333 161535 9336
rect 161477 9327 161535 9333
rect 168377 9333 168389 9336
rect 168423 9333 168435 9367
rect 168668 9364 168696 9404
rect 169588 9404 176654 9432
rect 169588 9364 169616 9404
rect 168668 9336 169616 9364
rect 170033 9367 170091 9373
rect 168377 9327 168435 9333
rect 170033 9333 170045 9367
rect 170079 9364 170091 9367
rect 170309 9367 170367 9373
rect 170309 9364 170321 9367
rect 170079 9336 170321 9364
rect 170079 9333 170091 9336
rect 170033 9327 170091 9333
rect 170309 9333 170321 9336
rect 170355 9333 170367 9367
rect 176626 9364 176654 9404
rect 185596 9404 186084 9432
rect 185489 9367 185547 9373
rect 185489 9364 185501 9367
rect 176626 9336 185501 9364
rect 170309 9327 170367 9333
rect 185489 9333 185501 9336
rect 185535 9333 185547 9367
rect 185489 9327 185547 9333
rect 185397 9299 185455 9305
rect 185397 9296 185409 9299
rect 157306 9268 161612 9296
rect 142203 9265 142215 9268
rect 142157 9259 142215 9265
rect 154025 9231 154083 9237
rect 154025 9197 154037 9231
rect 154071 9228 154083 9231
rect 161477 9231 161535 9237
rect 161477 9228 161489 9231
rect 154071 9200 161489 9228
rect 154071 9197 154083 9200
rect 154025 9191 154083 9197
rect 161477 9197 161489 9200
rect 161523 9197 161535 9231
rect 161477 9191 161535 9197
rect 35713 9163 35771 9169
rect 35713 9129 35725 9163
rect 35759 9160 35771 9163
rect 161584 9160 161612 9268
rect 170324 9268 185409 9296
rect 170324 9240 170352 9268
rect 185397 9265 185409 9268
rect 185443 9265 185455 9299
rect 185397 9259 185455 9265
rect 168469 9231 168527 9237
rect 168469 9228 168481 9231
rect 164206 9200 168481 9228
rect 164206 9160 164234 9200
rect 168469 9197 168481 9200
rect 168515 9197 168527 9231
rect 168469 9191 168527 9197
rect 170306 9188 170312 9240
rect 170364 9188 170370 9240
rect 171781 9231 171839 9237
rect 171781 9197 171793 9231
rect 171827 9228 171839 9231
rect 185596 9228 185624 9404
rect 185762 9364 185768 9376
rect 185723 9336 185768 9364
rect 185762 9324 185768 9336
rect 185820 9324 185826 9376
rect 171827 9200 185624 9228
rect 186056 9228 186084 9404
rect 233881 9401 233893 9435
rect 233927 9432 233939 9435
rect 243449 9435 243507 9441
rect 243449 9432 243461 9435
rect 233927 9404 243461 9432
rect 233927 9401 233939 9404
rect 233881 9395 233939 9401
rect 243449 9401 243461 9404
rect 243495 9401 243507 9435
rect 243556 9432 243584 9472
rect 244274 9460 244280 9472
rect 244332 9460 244338 9512
rect 244384 9509 244412 9540
rect 244550 9528 244556 9540
rect 244608 9528 244614 9580
rect 244642 9528 244648 9580
rect 244700 9568 244706 9580
rect 244829 9571 244887 9577
rect 244700 9540 244745 9568
rect 244700 9528 244706 9540
rect 244829 9537 244841 9571
rect 244875 9568 244887 9571
rect 245565 9571 245623 9577
rect 245565 9568 245577 9571
rect 244875 9540 245577 9568
rect 244875 9537 244887 9540
rect 244829 9531 244887 9537
rect 245565 9537 245577 9540
rect 245611 9537 245623 9571
rect 245565 9531 245623 9537
rect 247865 9571 247923 9577
rect 247865 9537 247877 9571
rect 247911 9568 247923 9571
rect 248233 9571 248291 9577
rect 248233 9568 248245 9571
rect 247911 9540 248245 9568
rect 247911 9537 247923 9540
rect 247865 9531 247923 9537
rect 248233 9537 248245 9540
rect 248279 9537 248291 9571
rect 270678 9568 270684 9580
rect 248233 9531 248291 9537
rect 253906 9540 270684 9568
rect 244369 9503 244427 9509
rect 244369 9469 244381 9503
rect 244415 9469 244427 9503
rect 253906 9500 253934 9540
rect 270678 9528 270684 9540
rect 270736 9528 270742 9580
rect 270862 9568 270868 9580
rect 270823 9540 270868 9568
rect 270862 9528 270868 9540
rect 270920 9528 270926 9580
rect 272328 9571 272386 9577
rect 272328 9537 272340 9571
rect 272374 9568 272386 9571
rect 272444 9568 272472 9646
rect 272374 9540 272472 9568
rect 272374 9537 272386 9540
rect 272328 9531 272386 9537
rect 273162 9528 273168 9580
rect 273220 9568 273226 9580
rect 273220 9566 277440 9568
rect 277504 9566 277532 9676
rect 277762 9664 277768 9676
rect 277820 9704 277826 9716
rect 278041 9707 278099 9713
rect 278041 9704 278053 9707
rect 277820 9676 278053 9704
rect 277820 9664 277826 9676
rect 278041 9673 278053 9676
rect 278087 9673 278099 9707
rect 278041 9667 278099 9673
rect 278130 9596 278136 9648
rect 278188 9636 278194 9648
rect 469398 9636 469404 9648
rect 278188 9608 469404 9636
rect 278188 9596 278194 9608
rect 469398 9596 469404 9608
rect 469456 9596 469462 9648
rect 273220 9540 277532 9566
rect 273220 9528 273226 9540
rect 277412 9538 277532 9540
rect 277670 9528 277676 9580
rect 277728 9568 277734 9580
rect 277857 9571 277915 9577
rect 277857 9568 277869 9571
rect 277728 9540 277869 9568
rect 277728 9528 277734 9540
rect 277857 9537 277869 9540
rect 277903 9568 277915 9571
rect 310698 9568 310704 9580
rect 277903 9540 310704 9568
rect 277903 9537 277915 9540
rect 277857 9531 277915 9537
rect 310698 9528 310704 9540
rect 310756 9528 310762 9580
rect 317322 9528 317328 9580
rect 317380 9568 317386 9580
rect 495434 9568 495440 9580
rect 317380 9540 495440 9568
rect 317380 9528 317386 9540
rect 495434 9528 495440 9540
rect 495492 9528 495498 9580
rect 244369 9463 244427 9469
rect 244476 9472 253934 9500
rect 258736 9472 261708 9500
rect 244476 9432 244504 9472
rect 245105 9435 245163 9441
rect 243556 9404 244504 9432
rect 244568 9404 244964 9432
rect 243449 9395 243507 9401
rect 191193 9367 191251 9373
rect 191193 9333 191205 9367
rect 191239 9364 191251 9367
rect 244568 9364 244596 9404
rect 191239 9336 244596 9364
rect 244936 9364 244964 9404
rect 245105 9401 245117 9435
rect 245151 9432 245163 9435
rect 258629 9435 258687 9441
rect 258629 9432 258641 9435
rect 245151 9404 258641 9432
rect 245151 9401 245163 9404
rect 245105 9395 245163 9401
rect 258629 9401 258641 9404
rect 258675 9401 258687 9435
rect 258629 9395 258687 9401
rect 258736 9364 258764 9472
rect 244936 9336 258764 9364
rect 258828 9404 261616 9432
rect 191239 9333 191251 9336
rect 191193 9327 191251 9333
rect 186225 9299 186283 9305
rect 186225 9265 186237 9299
rect 186271 9296 186283 9299
rect 258828 9296 258856 9404
rect 258905 9367 258963 9373
rect 258905 9333 258917 9367
rect 258951 9364 258963 9367
rect 261294 9364 261300 9376
rect 258951 9336 261300 9364
rect 258951 9333 258963 9336
rect 258905 9327 258963 9333
rect 261294 9324 261300 9336
rect 261352 9324 261358 9376
rect 261478 9364 261484 9376
rect 261439 9336 261484 9364
rect 261478 9324 261484 9336
rect 261536 9324 261542 9376
rect 186271 9268 238754 9296
rect 186271 9265 186283 9268
rect 186225 9259 186283 9265
rect 233881 9231 233939 9237
rect 233881 9228 233893 9231
rect 186056 9200 233893 9228
rect 171827 9197 171839 9200
rect 171781 9191 171839 9197
rect 233881 9197 233893 9200
rect 233927 9197 233939 9231
rect 233881 9191 233939 9197
rect 170122 9160 170128 9172
rect 35759 9132 161474 9160
rect 161584 9132 164234 9160
rect 168392 9132 170128 9160
rect 35759 9129 35771 9132
rect 35713 9123 35771 9129
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 150345 9095 150403 9101
rect 150345 9092 150357 9095
rect 7892 9064 150357 9092
rect 7892 9052 7898 9064
rect 150345 9061 150357 9064
rect 150391 9061 150403 9095
rect 150345 9055 150403 9061
rect 150529 9095 150587 9101
rect 150529 9061 150541 9095
rect 150575 9092 150587 9095
rect 154025 9095 154083 9101
rect 154025 9092 154037 9095
rect 150575 9064 154037 9092
rect 150575 9061 150587 9064
rect 150529 9055 150587 9061
rect 154025 9061 154037 9064
rect 154071 9061 154083 9095
rect 161446 9092 161474 9132
rect 168392 9092 168420 9132
rect 170122 9120 170128 9132
rect 170180 9120 170186 9172
rect 170398 9120 170404 9172
rect 170456 9160 170462 9172
rect 238726 9160 238754 9268
rect 248386 9268 258856 9296
rect 261588 9296 261616 9404
rect 261680 9364 261708 9472
rect 261754 9460 261760 9512
rect 261812 9500 261818 9512
rect 266817 9503 266875 9509
rect 266817 9500 266829 9503
rect 261812 9472 266829 9500
rect 261812 9460 261818 9472
rect 266817 9469 266829 9472
rect 266863 9469 266875 9503
rect 270954 9500 270960 9512
rect 266817 9463 266875 9469
rect 267016 9472 270960 9500
rect 267016 9364 267044 9472
rect 270954 9460 270960 9472
rect 271012 9460 271018 9512
rect 271049 9503 271107 9509
rect 271049 9469 271061 9503
rect 271095 9469 271107 9503
rect 271417 9503 271475 9509
rect 271417 9500 271429 9503
rect 271049 9463 271107 9469
rect 271248 9472 271429 9500
rect 267093 9435 267151 9441
rect 267093 9401 267105 9435
rect 267139 9432 267151 9435
rect 271064 9432 271092 9463
rect 271248 9432 271276 9472
rect 271417 9469 271429 9472
rect 271463 9469 271475 9503
rect 272058 9500 272064 9512
rect 271971 9472 272064 9500
rect 271417 9463 271475 9469
rect 272058 9460 272064 9472
rect 272116 9460 272122 9512
rect 277581 9503 277639 9509
rect 277581 9469 277593 9503
rect 277627 9500 277639 9503
rect 282181 9503 282239 9509
rect 282181 9500 282193 9503
rect 277627 9472 282193 9500
rect 277627 9469 277639 9472
rect 277581 9463 277639 9469
rect 282181 9469 282193 9472
rect 282227 9469 282239 9503
rect 282181 9463 282239 9469
rect 282273 9503 282331 9509
rect 282273 9469 282285 9503
rect 282319 9500 282331 9503
rect 445754 9500 445760 9512
rect 282319 9472 445760 9500
rect 282319 9469 282331 9472
rect 282273 9463 282331 9469
rect 445754 9460 445760 9472
rect 445812 9460 445818 9512
rect 267139 9404 270632 9432
rect 271064 9404 271276 9432
rect 267139 9401 267151 9404
rect 267093 9395 267151 9401
rect 261680 9336 267044 9364
rect 267185 9367 267243 9373
rect 267185 9333 267197 9367
rect 267231 9364 267243 9367
rect 270497 9367 270555 9373
rect 270497 9364 270509 9367
rect 267231 9336 270509 9364
rect 267231 9333 267243 9336
rect 267185 9327 267243 9333
rect 270497 9333 270509 9336
rect 270543 9333 270555 9367
rect 270604 9364 270632 9404
rect 271322 9392 271328 9444
rect 271380 9432 271386 9444
rect 272076 9432 272104 9460
rect 496354 9432 496360 9444
rect 271380 9404 272104 9432
rect 273226 9404 496360 9432
rect 271380 9392 271386 9404
rect 273226 9364 273254 9404
rect 496354 9392 496360 9404
rect 496412 9392 496418 9444
rect 273438 9364 273444 9376
rect 270604 9336 273254 9364
rect 273399 9336 273444 9364
rect 270497 9327 270555 9333
rect 273438 9324 273444 9336
rect 273496 9364 273502 9376
rect 273717 9367 273775 9373
rect 273496 9336 273668 9364
rect 273496 9324 273502 9336
rect 261588 9268 263916 9296
rect 248386 9160 248414 9268
rect 253293 9231 253351 9237
rect 253293 9197 253305 9231
rect 253339 9228 253351 9231
rect 253339 9200 258856 9228
rect 253339 9197 253351 9200
rect 253293 9191 253351 9197
rect 258828 9160 258856 9200
rect 261588 9200 263824 9228
rect 261588 9160 261616 9200
rect 263597 9163 263655 9169
rect 263597 9160 263609 9163
rect 170456 9132 233924 9160
rect 238726 9132 248414 9160
rect 248616 9132 258764 9160
rect 258828 9132 261616 9160
rect 261680 9132 263609 9160
rect 170456 9120 170462 9132
rect 161446 9064 168420 9092
rect 168469 9095 168527 9101
rect 154025 9055 154083 9061
rect 168469 9061 168481 9095
rect 168515 9092 168527 9095
rect 170214 9092 170220 9104
rect 168515 9064 170220 9092
rect 168515 9061 168527 9064
rect 168469 9055 168527 9061
rect 170214 9052 170220 9064
rect 170272 9052 170278 9104
rect 170309 9095 170367 9101
rect 170309 9061 170321 9095
rect 170355 9092 170367 9095
rect 233789 9095 233847 9101
rect 233789 9092 233801 9095
rect 170355 9064 233801 9092
rect 170355 9061 170367 9064
rect 170309 9055 170367 9061
rect 233789 9061 233801 9064
rect 233835 9061 233847 9095
rect 233896 9092 233924 9132
rect 248616 9092 248644 9132
rect 233896 9064 248644 9092
rect 253109 9095 253167 9101
rect 233789 9055 233847 9061
rect 253109 9061 253121 9095
rect 253155 9092 253167 9095
rect 258629 9095 258687 9101
rect 258629 9092 258641 9095
rect 253155 9064 258641 9092
rect 253155 9061 253167 9064
rect 253109 9055 253167 9061
rect 258629 9061 258641 9064
rect 258675 9061 258687 9095
rect 258736 9092 258764 9132
rect 261680 9092 261708 9132
rect 263597 9129 263609 9132
rect 263643 9129 263655 9163
rect 263597 9123 263655 9129
rect 258736 9064 261708 9092
rect 261757 9095 261815 9101
rect 258629 9055 258687 9061
rect 261757 9061 261769 9095
rect 261803 9092 261815 9095
rect 263689 9095 263747 9101
rect 263689 9092 263701 9095
rect 261803 9064 263701 9092
rect 261803 9061 261815 9064
rect 261757 9055 261815 9061
rect 263689 9061 263701 9064
rect 263735 9061 263747 9095
rect 263796 9092 263824 9200
rect 263888 9160 263916 9268
rect 273640 9228 273668 9336
rect 273717 9333 273729 9367
rect 273763 9364 273775 9367
rect 277486 9364 277492 9376
rect 273763 9336 277492 9364
rect 273763 9333 273775 9336
rect 273717 9327 273775 9333
rect 277486 9324 277492 9336
rect 277544 9324 277550 9376
rect 277578 9324 277584 9376
rect 277636 9364 277642 9376
rect 455414 9364 455420 9376
rect 277636 9336 455420 9364
rect 277636 9324 277642 9336
rect 455414 9324 455420 9336
rect 455472 9324 455478 9376
rect 278133 9299 278191 9305
rect 278133 9265 278145 9299
rect 278179 9296 278191 9299
rect 280801 9299 280859 9305
rect 280801 9296 280813 9299
rect 278179 9268 280813 9296
rect 278179 9265 278191 9268
rect 278133 9259 278191 9265
rect 280801 9265 280813 9268
rect 280847 9265 280859 9299
rect 280801 9259 280859 9265
rect 280890 9256 280896 9308
rect 280948 9296 280954 9308
rect 382550 9296 382556 9308
rect 280948 9268 382556 9296
rect 280948 9256 280954 9268
rect 382550 9256 382556 9268
rect 382608 9256 382614 9308
rect 273640 9200 277624 9228
rect 277596 9160 277624 9200
rect 278038 9188 278044 9240
rect 278096 9228 278102 9240
rect 282089 9231 282147 9237
rect 282089 9228 282101 9231
rect 278096 9200 282101 9228
rect 278096 9188 278102 9200
rect 282089 9197 282101 9200
rect 282135 9197 282147 9231
rect 282089 9191 282147 9197
rect 282181 9231 282239 9237
rect 282181 9197 282193 9231
rect 282227 9228 282239 9231
rect 360102 9228 360108 9240
rect 282227 9200 360108 9228
rect 282227 9197 282239 9200
rect 282181 9191 282239 9197
rect 360102 9188 360108 9200
rect 360160 9188 360166 9240
rect 469674 9160 469680 9172
rect 263888 9132 277532 9160
rect 277596 9132 469680 9160
rect 277397 9095 277455 9101
rect 277397 9092 277409 9095
rect 263796 9064 277409 9092
rect 263689 9055 263747 9061
rect 277397 9061 277409 9064
rect 277443 9061 277455 9095
rect 277504 9092 277532 9132
rect 469674 9120 469680 9132
rect 469732 9120 469738 9172
rect 280890 9092 280896 9104
rect 277504 9064 280896 9092
rect 277397 9055 277455 9061
rect 280890 9052 280896 9064
rect 280948 9052 280954 9104
rect 280985 9095 281043 9101
rect 280985 9061 280997 9095
rect 281031 9092 281043 9095
rect 282086 9092 282092 9104
rect 281031 9064 282092 9092
rect 281031 9061 281043 9064
rect 280985 9055 281043 9061
rect 282086 9052 282092 9064
rect 282144 9052 282150 9104
rect 282181 9095 282239 9101
rect 282181 9061 282193 9095
rect 282227 9092 282239 9095
rect 401226 9092 401232 9104
rect 282227 9064 401232 9092
rect 282227 9061 282239 9064
rect 282181 9055 282239 9061
rect 401226 9052 401232 9064
rect 401284 9052 401290 9104
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 138385 9027 138443 9033
rect 138385 9024 138397 9027
rect 4028 8996 138397 9024
rect 4028 8984 4034 8996
rect 138385 8993 138397 8996
rect 138431 8993 138443 9027
rect 138385 8987 138443 8993
rect 147766 8984 147772 9036
rect 147824 9024 147830 9036
rect 372982 9024 372988 9036
rect 147824 8996 372988 9024
rect 147824 8984 147830 8996
rect 372982 8984 372988 8996
rect 373040 8984 373046 9036
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 115937 8959 115995 8965
rect 115937 8956 115949 8959
rect 9272 8928 115949 8956
rect 9272 8916 9278 8928
rect 115937 8925 115949 8928
rect 115983 8925 115995 8959
rect 115937 8919 115995 8925
rect 116578 8916 116584 8968
rect 116636 8956 116642 8968
rect 117038 8956 117044 8968
rect 116636 8928 117044 8956
rect 116636 8916 116642 8928
rect 117038 8916 117044 8928
rect 117096 8956 117102 8968
rect 341150 8956 341156 8968
rect 117096 8928 147674 8956
rect 117096 8916 117102 8928
rect 147646 8888 147674 8928
rect 147784 8928 341156 8956
rect 147784 8888 147812 8928
rect 341150 8916 341156 8928
rect 341208 8916 341214 8968
rect 147646 8860 147812 8888
rect 150345 8891 150403 8897
rect 150345 8857 150357 8891
rect 150391 8888 150403 8891
rect 150986 8888 150992 8900
rect 150391 8860 150992 8888
rect 150391 8857 150403 8860
rect 150345 8851 150403 8857
rect 150986 8848 150992 8860
rect 151044 8888 151050 8900
rect 153013 8891 153071 8897
rect 153013 8888 153025 8891
rect 151044 8860 153025 8888
rect 151044 8848 151050 8860
rect 153013 8857 153025 8860
rect 153059 8857 153071 8891
rect 153013 8851 153071 8857
rect 153105 8891 153163 8897
rect 153105 8857 153117 8891
rect 153151 8888 153163 8891
rect 241517 8891 241575 8897
rect 241517 8888 241529 8891
rect 153151 8860 241529 8888
rect 153151 8857 153163 8860
rect 153105 8851 153163 8857
rect 241517 8857 241529 8860
rect 241563 8857 241575 8891
rect 241517 8851 241575 8857
rect 243449 8891 243507 8897
rect 243449 8857 243461 8891
rect 243495 8888 243507 8891
rect 253293 8891 253351 8897
rect 253293 8888 253305 8891
rect 243495 8860 253305 8888
rect 243495 8857 243507 8860
rect 243449 8851 243507 8857
rect 253293 8857 253305 8860
rect 253339 8857 253351 8891
rect 253293 8851 253351 8857
rect 253385 8891 253443 8897
rect 253385 8857 253397 8891
rect 253431 8888 253443 8891
rect 451458 8888 451464 8900
rect 253431 8860 451464 8888
rect 253431 8857 253443 8860
rect 253385 8851 253443 8857
rect 451458 8848 451464 8860
rect 451516 8848 451522 8900
rect 116029 8823 116087 8829
rect 116029 8789 116041 8823
rect 116075 8820 116087 8823
rect 230385 8823 230443 8829
rect 230385 8820 230397 8823
rect 116075 8792 230397 8820
rect 116075 8789 116087 8792
rect 116029 8783 116087 8789
rect 230385 8789 230397 8792
rect 230431 8789 230443 8823
rect 230385 8783 230443 8789
rect 233789 8823 233847 8829
rect 233789 8789 233801 8823
rect 233835 8820 233847 8823
rect 253109 8823 253167 8829
rect 253109 8820 253121 8823
rect 233835 8792 253121 8820
rect 233835 8789 233847 8792
rect 233789 8783 233847 8789
rect 253109 8789 253121 8792
rect 253155 8789 253167 8823
rect 253109 8783 253167 8789
rect 253201 8823 253259 8829
rect 253201 8789 253213 8823
rect 253247 8820 253259 8823
rect 258537 8823 258595 8829
rect 258537 8820 258549 8823
rect 253247 8792 258549 8820
rect 253247 8789 253259 8792
rect 253201 8783 253259 8789
rect 258537 8789 258549 8792
rect 258583 8789 258595 8823
rect 258537 8783 258595 8789
rect 258629 8823 258687 8829
rect 258629 8789 258641 8823
rect 258675 8820 258687 8823
rect 261665 8823 261723 8829
rect 261665 8820 261677 8823
rect 258675 8792 261677 8820
rect 258675 8789 258687 8792
rect 258629 8783 258687 8789
rect 261665 8789 261677 8792
rect 261711 8789 261723 8823
rect 261665 8783 261723 8789
rect 261757 8823 261815 8829
rect 261757 8789 261769 8823
rect 261803 8820 261815 8823
rect 268381 8823 268439 8829
rect 261803 8792 267688 8820
rect 261803 8789 261815 8792
rect 261757 8783 261815 8789
rect 3878 8712 3884 8764
rect 3936 8752 3942 8764
rect 120077 8755 120135 8761
rect 120077 8752 120089 8755
rect 3936 8724 120089 8752
rect 3936 8712 3942 8724
rect 120077 8721 120089 8724
rect 120123 8721 120135 8755
rect 120077 8715 120135 8721
rect 148965 8755 149023 8761
rect 148965 8721 148977 8755
rect 149011 8752 149023 8755
rect 267185 8755 267243 8761
rect 267185 8752 267197 8755
rect 149011 8724 267197 8752
rect 149011 8721 149023 8724
rect 148965 8715 149023 8721
rect 267185 8721 267197 8724
rect 267231 8721 267243 8755
rect 267660 8752 267688 8792
rect 268381 8789 268393 8823
rect 268427 8820 268439 8823
rect 279329 8823 279387 8829
rect 268427 8792 279280 8820
rect 268427 8789 268439 8792
rect 268381 8783 268439 8789
rect 279145 8755 279203 8761
rect 279145 8752 279157 8755
rect 267660 8724 279157 8752
rect 267185 8715 267243 8721
rect 279145 8721 279157 8724
rect 279191 8721 279203 8755
rect 279252 8752 279280 8792
rect 279329 8789 279341 8823
rect 279375 8820 279387 8823
rect 321462 8820 321468 8832
rect 279375 8792 321468 8820
rect 279375 8789 279387 8792
rect 279329 8783 279387 8789
rect 321462 8780 321468 8792
rect 321520 8780 321526 8832
rect 282181 8755 282239 8761
rect 282181 8752 282193 8755
rect 279252 8724 282193 8752
rect 279145 8715 279203 8721
rect 282181 8721 282193 8724
rect 282227 8721 282239 8755
rect 282181 8715 282239 8721
rect 282273 8755 282331 8761
rect 282273 8721 282285 8755
rect 282319 8752 282331 8755
rect 467742 8752 467748 8764
rect 282319 8724 467748 8752
rect 282319 8721 282331 8724
rect 282273 8715 282331 8721
rect 467742 8712 467748 8724
rect 467800 8712 467806 8764
rect 6730 8644 6736 8696
rect 6788 8684 6794 8696
rect 150437 8687 150495 8693
rect 150437 8684 150449 8687
rect 6788 8656 150449 8684
rect 6788 8644 6794 8656
rect 150437 8653 150449 8656
rect 150483 8653 150495 8687
rect 150437 8647 150495 8653
rect 152921 8687 152979 8693
rect 152921 8653 152933 8687
rect 152967 8684 152979 8687
rect 320450 8684 320456 8696
rect 152967 8656 320456 8684
rect 152967 8653 152979 8656
rect 152921 8647 152979 8653
rect 320450 8644 320456 8656
rect 320508 8644 320514 8696
rect 77481 8619 77539 8625
rect 77481 8585 77493 8619
rect 77527 8616 77539 8619
rect 168285 8619 168343 8625
rect 168285 8616 168297 8619
rect 77527 8588 168297 8616
rect 77527 8585 77539 8588
rect 77481 8579 77539 8585
rect 168285 8585 168297 8588
rect 168331 8585 168343 8619
rect 168285 8579 168343 8585
rect 168377 8619 168435 8625
rect 168377 8585 168389 8619
rect 168423 8616 168435 8619
rect 171781 8619 171839 8625
rect 171781 8616 171793 8619
rect 168423 8588 171793 8616
rect 168423 8585 168435 8588
rect 168377 8579 168435 8585
rect 171781 8585 171793 8588
rect 171827 8585 171839 8619
rect 171781 8579 171839 8585
rect 230385 8619 230443 8625
rect 230385 8585 230397 8619
rect 230431 8616 230443 8619
rect 253201 8619 253259 8625
rect 253201 8616 253213 8619
rect 230431 8588 253213 8616
rect 230431 8585 230443 8588
rect 230385 8579 230443 8585
rect 253201 8585 253213 8588
rect 253247 8585 253259 8619
rect 253201 8579 253259 8585
rect 258537 8619 258595 8625
rect 258537 8585 258549 8619
rect 258583 8616 258595 8619
rect 261757 8619 261815 8625
rect 261757 8616 261769 8619
rect 258583 8588 261769 8616
rect 258583 8585 258595 8588
rect 258537 8579 258595 8585
rect 261757 8585 261769 8588
rect 261803 8585 261815 8619
rect 261757 8579 261815 8585
rect 263689 8619 263747 8625
rect 263689 8585 263701 8619
rect 263735 8616 263747 8619
rect 268381 8619 268439 8625
rect 268381 8616 268393 8619
rect 263735 8588 268393 8616
rect 263735 8585 263747 8588
rect 263689 8579 263747 8585
rect 268381 8585 268393 8588
rect 268427 8585 268439 8619
rect 273717 8619 273775 8625
rect 273717 8616 273729 8619
rect 268381 8579 268439 8585
rect 268488 8588 273729 8616
rect 76745 8551 76803 8557
rect 76745 8517 76757 8551
rect 76791 8548 76803 8551
rect 168466 8548 168472 8560
rect 76791 8520 168472 8548
rect 76791 8517 76803 8520
rect 76745 8511 76803 8517
rect 168466 8508 168472 8520
rect 168524 8508 168530 8560
rect 168650 8508 168656 8560
rect 168708 8548 168714 8560
rect 263781 8551 263839 8557
rect 168708 8520 263732 8548
rect 168708 8508 168714 8520
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 4948 8452 238754 8480
rect 4948 8440 4954 8452
rect 7006 8372 7012 8424
rect 7064 8412 7070 8424
rect 148505 8415 148563 8421
rect 148505 8412 148517 8415
rect 7064 8384 148517 8412
rect 7064 8372 7070 8384
rect 148505 8381 148517 8384
rect 148551 8412 148563 8415
rect 153105 8415 153163 8421
rect 153105 8412 153117 8415
rect 148551 8384 153117 8412
rect 148551 8381 148563 8384
rect 148505 8375 148563 8381
rect 153105 8381 153117 8384
rect 153151 8381 153163 8415
rect 153105 8375 153163 8381
rect 168285 8415 168343 8421
rect 168285 8381 168297 8415
rect 168331 8412 168343 8415
rect 170309 8415 170367 8421
rect 170309 8412 170321 8415
rect 168331 8384 170321 8412
rect 168331 8381 168343 8384
rect 168285 8375 168343 8381
rect 170309 8381 170321 8384
rect 170355 8381 170367 8415
rect 238726 8412 238754 8452
rect 240042 8440 240048 8492
rect 240100 8480 240106 8492
rect 245105 8483 245163 8489
rect 245105 8480 245117 8483
rect 240100 8452 245117 8480
rect 240100 8440 240106 8452
rect 245105 8449 245117 8452
rect 245151 8449 245163 8483
rect 245105 8443 245163 8449
rect 245565 8483 245623 8489
rect 245565 8449 245577 8483
rect 245611 8480 245623 8483
rect 253385 8483 253443 8489
rect 253385 8480 253397 8483
rect 245611 8452 253397 8480
rect 245611 8449 245623 8452
rect 245565 8443 245623 8449
rect 253385 8449 253397 8452
rect 253431 8449 253443 8483
rect 263597 8483 263655 8489
rect 263597 8480 263609 8483
rect 253385 8443 253443 8449
rect 253906 8452 263609 8480
rect 244642 8412 244648 8424
rect 238726 8384 244648 8412
rect 170309 8375 170367 8381
rect 244642 8372 244648 8384
rect 244700 8372 244706 8424
rect 247865 8415 247923 8421
rect 247865 8381 247877 8415
rect 247911 8412 247923 8415
rect 253906 8412 253934 8452
rect 263597 8449 263609 8452
rect 263643 8449 263655 8483
rect 263597 8443 263655 8449
rect 247911 8384 253934 8412
rect 263704 8412 263732 8520
rect 263781 8517 263793 8551
rect 263827 8548 263839 8551
rect 268488 8548 268516 8588
rect 273717 8585 273729 8588
rect 273763 8585 273775 8619
rect 273717 8579 273775 8585
rect 273806 8576 273812 8628
rect 273864 8616 273870 8628
rect 277670 8616 277676 8628
rect 273864 8588 277676 8616
rect 273864 8576 273870 8588
rect 277670 8576 277676 8588
rect 277728 8576 277734 8628
rect 277765 8619 277823 8625
rect 277765 8585 277777 8619
rect 277811 8616 277823 8619
rect 405366 8616 405372 8628
rect 277811 8588 405372 8616
rect 277811 8585 277823 8588
rect 277765 8579 277823 8585
rect 405366 8576 405372 8588
rect 405424 8576 405430 8628
rect 263827 8520 268516 8548
rect 271417 8551 271475 8557
rect 263827 8517 263839 8520
rect 263781 8511 263839 8517
rect 271417 8517 271429 8551
rect 271463 8548 271475 8551
rect 282181 8551 282239 8557
rect 282181 8548 282193 8551
rect 271463 8520 282193 8548
rect 271463 8517 271475 8520
rect 271417 8511 271475 8517
rect 282181 8517 282193 8520
rect 282227 8517 282239 8551
rect 282181 8511 282239 8517
rect 282270 8508 282276 8560
rect 282328 8548 282334 8560
rect 343910 8548 343916 8560
rect 282328 8520 343916 8548
rect 282328 8508 282334 8520
rect 343910 8508 343916 8520
rect 343968 8508 343974 8560
rect 263873 8483 263931 8489
rect 263873 8449 263885 8483
rect 263919 8480 263931 8483
rect 340874 8480 340880 8492
rect 263919 8452 340880 8480
rect 263919 8449 263931 8452
rect 263873 8443 263931 8449
rect 340874 8440 340880 8452
rect 340932 8440 340938 8492
rect 271322 8412 271328 8424
rect 263704 8384 271328 8412
rect 247911 8381 247923 8384
rect 247865 8375 247923 8381
rect 271322 8372 271328 8384
rect 271380 8372 271386 8424
rect 271509 8415 271567 8421
rect 271509 8381 271521 8415
rect 271555 8412 271567 8415
rect 277765 8415 277823 8421
rect 277765 8412 277777 8415
rect 271555 8384 277777 8412
rect 271555 8381 271567 8384
rect 271509 8375 271567 8381
rect 277765 8381 277777 8384
rect 277811 8381 277823 8415
rect 277765 8375 277823 8381
rect 278041 8415 278099 8421
rect 278041 8381 278053 8415
rect 278087 8412 278099 8415
rect 282089 8415 282147 8421
rect 282089 8412 282101 8415
rect 278087 8384 282101 8412
rect 278087 8381 278099 8384
rect 278041 8375 278099 8381
rect 282089 8381 282101 8384
rect 282135 8381 282147 8415
rect 282089 8375 282147 8381
rect 282181 8415 282239 8421
rect 282181 8381 282193 8415
rect 282227 8412 282239 8415
rect 328270 8412 328276 8424
rect 282227 8384 328276 8412
rect 282227 8381 282239 8384
rect 282181 8375 282239 8381
rect 328270 8372 328276 8384
rect 328328 8372 328334 8424
rect 66165 8347 66223 8353
rect 66165 8313 66177 8347
rect 66211 8344 66223 8347
rect 468018 8344 468024 8356
rect 66211 8316 468024 8344
rect 66211 8313 66223 8316
rect 66165 8307 66223 8313
rect 468018 8304 468024 8316
rect 468076 8304 468082 8356
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 16666 8276 16672 8288
rect 5500 8248 16672 8276
rect 5500 8236 5506 8248
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 301498 8236 301504 8288
rect 301556 8276 301562 8288
rect 310974 8276 310980 8288
rect 301556 8248 310980 8276
rect 301556 8236 301562 8248
rect 310974 8236 310980 8248
rect 311032 8236 311038 8288
rect 8570 8168 8576 8220
rect 8628 8208 8634 8220
rect 23290 8208 23296 8220
rect 8628 8180 23296 8208
rect 8628 8168 8634 8180
rect 23290 8168 23296 8180
rect 23348 8168 23354 8220
rect 308122 8168 308128 8220
rect 308180 8208 308186 8220
rect 404998 8208 405004 8220
rect 308180 8180 405004 8208
rect 308180 8168 308186 8180
rect 404998 8168 405004 8180
rect 405056 8168 405062 8220
rect 9582 8100 9588 8152
rect 9640 8140 9646 8152
rect 129274 8140 129280 8152
rect 9640 8112 129280 8140
rect 9640 8100 9646 8112
rect 129274 8100 129280 8112
rect 129332 8100 129338 8152
rect 222010 8100 222016 8152
rect 222068 8140 222074 8152
rect 444098 8140 444104 8152
rect 222068 8112 444104 8140
rect 222068 8100 222074 8112
rect 444098 8100 444104 8112
rect 444156 8100 444162 8152
rect 149146 8032 149152 8084
rect 149204 8072 149210 8084
rect 340414 8072 340420 8084
rect 149204 8044 340420 8072
rect 149204 8032 149210 8044
rect 340414 8032 340420 8044
rect 340472 8032 340478 8084
rect 42334 7964 42340 8016
rect 42392 8004 42398 8016
rect 215386 8004 215392 8016
rect 42392 7976 215392 8004
rect 42392 7964 42398 7976
rect 215386 7964 215392 7976
rect 215444 7964 215450 8016
rect 135898 7896 135904 7948
rect 135956 7936 135962 7948
rect 333054 7936 333060 7948
rect 135956 7908 333060 7936
rect 135956 7896 135962 7908
rect 333054 7896 333060 7908
rect 333112 7896 333118 7948
rect 88518 7828 88524 7880
rect 88576 7868 88582 7880
rect 89530 7868 89536 7880
rect 88576 7840 89536 7868
rect 88576 7828 88582 7840
rect 89530 7828 89536 7840
rect 89588 7868 89594 7880
rect 168650 7868 168656 7880
rect 89588 7840 168656 7868
rect 89588 7828 89594 7840
rect 168650 7828 168656 7840
rect 168708 7828 168714 7880
rect 203061 7871 203119 7877
rect 203061 7837 203073 7871
rect 203107 7868 203119 7871
rect 389818 7868 389824 7880
rect 203107 7840 389824 7868
rect 203107 7837 203119 7840
rect 203061 7831 203119 7837
rect 389818 7828 389824 7840
rect 389876 7828 389882 7880
rect 63034 7760 63040 7812
rect 63092 7800 63098 7812
rect 278590 7800 278596 7812
rect 63092 7772 278596 7800
rect 63092 7760 63098 7772
rect 278590 7760 278596 7772
rect 278648 7760 278654 7812
rect 36538 7692 36544 7744
rect 36596 7732 36602 7744
rect 272518 7732 272524 7744
rect 36596 7704 272524 7732
rect 36596 7692 36602 7704
rect 272518 7692 272524 7704
rect 272576 7692 272582 7744
rect 29914 7624 29920 7676
rect 29972 7664 29978 7676
rect 78582 7664 78588 7676
rect 29972 7636 78588 7664
rect 29972 7624 29978 7636
rect 78582 7624 78588 7636
rect 78640 7624 78646 7676
rect 23290 7556 23296 7608
rect 23348 7596 23354 7608
rect 75638 7596 75644 7608
rect 23348 7568 75644 7596
rect 23348 7556 23354 7568
rect 75638 7556 75644 7568
rect 75696 7556 75702 7608
rect 241882 7556 241888 7608
rect 241940 7596 241946 7608
rect 384574 7596 384580 7608
rect 241940 7568 384580 7596
rect 241940 7556 241946 7568
rect 384574 7556 384580 7568
rect 384632 7556 384638 7608
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 418338 7528 418344 7540
rect 10100 7500 418344 7528
rect 10100 7488 10106 7500
rect 418338 7488 418344 7500
rect 418396 7488 418402 7540
rect 69658 7420 69664 7472
rect 69716 7460 69722 7472
rect 310238 7460 310244 7472
rect 69716 7432 310244 7460
rect 69716 7420 69722 7432
rect 310238 7420 310244 7432
rect 310296 7420 310302 7472
rect 54478 5312 54484 5364
rect 54536 5352 54542 5364
rect 326522 5352 326528 5364
rect 54536 5324 326528 5352
rect 54536 5312 54542 5324
rect 326522 5312 326528 5324
rect 326580 5312 326586 5364
rect 60550 5244 60556 5296
rect 60608 5284 60614 5296
rect 342438 5284 342444 5296
rect 60608 5256 342444 5284
rect 60608 5244 60614 5256
rect 342438 5244 342444 5256
rect 342496 5244 342502 5296
rect 69100 5219 69158 5225
rect 69100 5185 69112 5219
rect 69146 5216 69158 5219
rect 318058 5216 318064 5228
rect 69146 5188 318064 5216
rect 69146 5185 69158 5188
rect 69100 5179 69158 5185
rect 318058 5176 318064 5188
rect 318116 5176 318122 5228
rect 8018 5108 8024 5160
rect 8076 5148 8082 5160
rect 68833 5151 68891 5157
rect 68833 5148 68845 5151
rect 8076 5120 68845 5148
rect 8076 5108 8082 5120
rect 68756 4808 68784 5120
rect 68833 5117 68845 5120
rect 68879 5117 68891 5151
rect 68833 5111 68891 5117
rect 205910 5040 205916 5092
rect 205968 5080 205974 5092
rect 376478 5080 376484 5092
rect 205968 5052 376484 5080
rect 205968 5040 205974 5052
rect 376478 5040 376484 5052
rect 376536 5040 376542 5092
rect 70213 5015 70271 5021
rect 70213 4981 70225 5015
rect 70259 5012 70271 5015
rect 339954 5012 339960 5024
rect 70259 4984 339960 5012
rect 70259 4981 70271 4984
rect 70213 4975 70271 4981
rect 339954 4972 339960 4984
rect 340012 4972 340018 5024
rect 88518 4808 88524 4820
rect 68756 4780 88524 4808
rect 88518 4768 88524 4780
rect 88576 4768 88582 4820
rect 148318 4768 148324 4820
rect 148376 4808 148382 4820
rect 470042 4808 470048 4820
rect 148376 4780 470048 4808
rect 148376 4768 148382 4780
rect 470042 4768 470048 4780
rect 470100 4768 470106 4820
rect 225509 4471 225567 4477
rect 225509 4437 225521 4471
rect 225555 4468 225567 4471
rect 349798 4468 349804 4480
rect 225555 4440 349804 4468
rect 225555 4437 225567 4440
rect 225509 4431 225567 4437
rect 349798 4428 349804 4440
rect 349856 4428 349862 4480
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 371234 4128 371240 4140
rect 9456 4100 371240 4128
rect 9456 4088 9462 4100
rect 371234 4088 371240 4100
rect 371292 4128 371298 4140
rect 372430 4128 372436 4140
rect 371292 4100 372436 4128
rect 371292 4088 371298 4100
rect 372430 4088 372436 4100
rect 372488 4088 372494 4140
rect 98822 4020 98828 4072
rect 98880 4060 98886 4072
rect 293678 4060 293684 4072
rect 98880 4032 293684 4060
rect 98880 4020 98886 4032
rect 293678 4020 293684 4032
rect 293736 4020 293742 4072
rect 302878 4020 302884 4072
rect 302936 4060 302942 4072
rect 310882 4060 310888 4072
rect 302936 4032 310888 4060
rect 302936 4020 302942 4032
rect 310882 4020 310888 4032
rect 310940 4020 310946 4072
rect 310977 4063 311035 4069
rect 310977 4029 310989 4063
rect 311023 4060 311035 4063
rect 315298 4060 315304 4072
rect 311023 4032 315304 4060
rect 311023 4029 311035 4032
rect 310977 4023 311035 4029
rect 315298 4020 315304 4032
rect 315356 4020 315362 4072
rect 318705 4063 318763 4069
rect 318705 4029 318717 4063
rect 318751 4060 318763 4063
rect 463326 4060 463332 4072
rect 318751 4032 463332 4060
rect 318751 4029 318763 4032
rect 318705 4023 318763 4029
rect 463326 4020 463332 4032
rect 463384 4020 463390 4072
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 193766 3992 193772 4004
rect 5040 3964 193772 3992
rect 5040 3952 5046 3964
rect 193766 3952 193772 3964
rect 193824 3952 193830 4004
rect 208854 3952 208860 4004
rect 208912 3992 208918 4004
rect 414842 3992 414848 4004
rect 208912 3964 414848 3992
rect 208912 3952 208918 3964
rect 414842 3952 414848 3964
rect 414900 3952 414906 4004
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 233142 3924 233148 3936
rect 9824 3896 233148 3924
rect 9824 3884 9830 3896
rect 233142 3884 233148 3896
rect 233200 3884 233206 3936
rect 434990 3924 434996 3936
rect 238726 3896 434996 3924
rect 8478 3816 8484 3868
rect 8536 3856 8542 3868
rect 236086 3856 236092 3868
rect 8536 3828 236092 3856
rect 8536 3816 8542 3828
rect 236086 3816 236092 3828
rect 236144 3856 236150 3868
rect 238726 3856 238754 3896
rect 434990 3884 434996 3896
rect 435048 3884 435054 3936
rect 236144 3828 238754 3856
rect 236144 3816 236150 3828
rect 257430 3816 257436 3868
rect 257488 3856 257494 3868
rect 493870 3856 493876 3868
rect 257488 3828 493876 3856
rect 257488 3816 257494 3828
rect 493870 3816 493876 3828
rect 493928 3816 493934 3868
rect 69566 3748 69572 3800
rect 69624 3788 69630 3800
rect 313826 3788 313832 3800
rect 69624 3760 313832 3788
rect 69624 3748 69630 3760
rect 313826 3748 313832 3760
rect 313884 3748 313890 3800
rect 315114 3748 315120 3800
rect 315172 3788 315178 3800
rect 475470 3788 475476 3800
rect 315172 3760 475476 3788
rect 315172 3748 315178 3760
rect 475470 3748 475476 3760
rect 475528 3748 475534 3800
rect 108942 3680 108948 3732
rect 109000 3720 109006 3732
rect 389358 3720 389364 3732
rect 109000 3692 389364 3720
rect 109000 3680 109006 3692
rect 389358 3680 389364 3692
rect 389416 3680 389422 3732
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 21174 3652 21180 3664
rect 8720 3624 21180 3652
rect 8720 3612 8726 3624
rect 21174 3612 21180 3624
rect 21232 3612 21238 3664
rect 39206 3612 39212 3664
rect 39264 3652 39270 3664
rect 338022 3652 338028 3664
rect 39264 3624 338028 3652
rect 39264 3612 39270 3624
rect 338022 3612 338028 3624
rect 338080 3612 338086 3664
rect 348326 3612 348332 3664
rect 348384 3652 348390 3664
rect 349062 3652 349068 3664
rect 348384 3624 349068 3652
rect 348384 3612 348390 3624
rect 349062 3612 349068 3624
rect 349120 3612 349126 3664
rect 360286 3612 360292 3664
rect 360344 3652 360350 3664
rect 361482 3652 361488 3664
rect 360344 3624 361488 3652
rect 360344 3612 360350 3624
rect 361482 3612 361488 3624
rect 361540 3612 361546 3664
rect 363414 3612 363420 3664
rect 363472 3652 363478 3664
rect 365806 3652 365812 3664
rect 363472 3624 365812 3652
rect 363472 3612 363478 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 369302 3612 369308 3664
rect 369360 3652 369366 3664
rect 460382 3652 460388 3664
rect 369360 3624 460388 3652
rect 369360 3612 369366 3624
rect 460382 3612 460388 3624
rect 460440 3612 460446 3664
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 24118 3584 24124 3596
rect 9916 3556 24124 3584
rect 9916 3544 9922 3556
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 63494 3544 63500 3596
rect 63552 3584 63558 3596
rect 376018 3584 376024 3596
rect 63552 3556 376024 3584
rect 63552 3544 63558 3556
rect 376018 3544 376024 3556
rect 376076 3544 376082 3596
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 33318 3516 33324 3528
rect 6052 3488 33324 3516
rect 6052 3476 6058 3488
rect 33318 3476 33324 3488
rect 33376 3476 33382 3528
rect 72234 3476 72240 3528
rect 72292 3516 72298 3528
rect 439038 3516 439044 3528
rect 72292 3488 439044 3516
rect 72292 3476 72298 3488
rect 439038 3476 439044 3488
rect 439096 3476 439102 3528
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 484486 3448 484492 3460
rect 8168 3420 484492 3448
rect 8168 3408 8174 3420
rect 484486 3408 484492 3420
rect 484544 3408 484550 3460
rect 14 3340 20 3392
rect 72 3380 78 3392
rect 117038 3380 117044 3392
rect 72 3352 117044 3380
rect 72 3340 78 3352
rect 117038 3340 117044 3352
rect 117096 3340 117102 3392
rect 145374 3340 145380 3392
rect 145432 3380 145438 3392
rect 310977 3383 311035 3389
rect 310977 3380 310989 3383
rect 145432 3352 310989 3380
rect 145432 3340 145438 3352
rect 310977 3349 310989 3352
rect 311023 3349 311035 3383
rect 310977 3343 311035 3349
rect 311250 3340 311256 3392
rect 311308 3380 311314 3392
rect 311894 3380 311900 3392
rect 311308 3352 311900 3380
rect 311308 3340 311314 3352
rect 311894 3340 311900 3352
rect 311952 3340 311958 3392
rect 312081 3383 312139 3389
rect 312081 3349 312093 3383
rect 312127 3380 312139 3383
rect 318705 3383 318763 3389
rect 318705 3380 318717 3383
rect 312127 3352 318717 3380
rect 312127 3349 312139 3352
rect 312081 3343 312139 3349
rect 318705 3349 318717 3352
rect 318751 3349 318763 3383
rect 318705 3343 318763 3349
rect 331858 3340 331864 3392
rect 331916 3380 331922 3392
rect 445110 3380 445116 3392
rect 331916 3352 445116 3380
rect 331916 3340 331922 3352
rect 445110 3340 445116 3352
rect 445168 3340 445174 3392
rect 157334 3272 157340 3324
rect 157392 3312 157398 3324
rect 311986 3312 311992 3324
rect 157392 3284 311992 3312
rect 157392 3272 157398 3284
rect 311986 3272 311992 3284
rect 312044 3272 312050 3324
rect 314378 3272 314384 3324
rect 314436 3312 314442 3324
rect 414934 3312 414940 3324
rect 314436 3284 414940 3312
rect 314436 3272 314442 3284
rect 414934 3272 414940 3284
rect 414992 3272 414998 3324
rect 172606 3204 172612 3256
rect 172664 3244 172670 3256
rect 322290 3244 322296 3256
rect 172664 3216 322296 3244
rect 172664 3204 172670 3216
rect 322290 3204 322296 3216
rect 322348 3204 322354 3256
rect 330478 3204 330484 3256
rect 330536 3244 330542 3256
rect 342254 3244 342260 3256
rect 330536 3216 342260 3244
rect 330536 3204 330542 3216
rect 342254 3204 342260 3216
rect 342312 3204 342318 3256
rect 366358 3204 366364 3256
rect 366416 3244 366422 3256
rect 436094 3244 436100 3256
rect 366416 3216 436100 3244
rect 366416 3204 366422 3216
rect 436094 3204 436100 3216
rect 436152 3204 436158 3256
rect 498197 3247 498255 3253
rect 498197 3213 498209 3247
rect 498243 3244 498255 3247
rect 499758 3244 499764 3256
rect 498243 3216 499764 3244
rect 498243 3213 498255 3216
rect 498197 3207 498255 3213
rect 499758 3204 499764 3216
rect 499816 3204 499822 3256
rect 45278 3136 45284 3188
rect 45336 3176 45342 3188
rect 182174 3176 182180 3188
rect 45336 3148 182180 3176
rect 45336 3136 45342 3148
rect 182174 3136 182180 3148
rect 182232 3136 182238 3188
rect 214926 3136 214932 3188
rect 214984 3176 214990 3188
rect 311342 3176 311348 3188
rect 214984 3148 311348 3176
rect 214984 3136 214990 3148
rect 311342 3136 311348 3148
rect 311400 3136 311406 3188
rect 311434 3136 311440 3188
rect 311492 3176 311498 3188
rect 454310 3176 454316 3188
rect 311492 3148 454316 3176
rect 311492 3136 311498 3148
rect 454310 3136 454316 3148
rect 454368 3136 454374 3188
rect 193766 3068 193772 3120
rect 193824 3108 193830 3120
rect 248414 3108 248420 3120
rect 193824 3080 248420 3108
rect 193824 3068 193830 3080
rect 248414 3068 248420 3080
rect 248472 3068 248478 3120
rect 287606 3068 287612 3120
rect 287664 3108 287670 3120
rect 420546 3108 420552 3120
rect 287664 3080 420552 3108
rect 287664 3068 287670 3080
rect 420546 3068 420552 3080
rect 420604 3068 420610 3120
rect 230198 3000 230204 3052
rect 230256 3040 230262 3052
rect 230256 3012 311112 3040
rect 230256 3000 230262 3012
rect 254302 2932 254308 2984
rect 254360 2972 254366 2984
rect 310514 2972 310520 2984
rect 254360 2944 310520 2972
rect 254360 2932 254366 2944
rect 310514 2932 310520 2944
rect 310572 2932 310578 2984
rect 311084 2972 311112 3012
rect 311158 3000 311164 3052
rect 311216 3040 311222 3052
rect 312081 3043 312139 3049
rect 312081 3040 312093 3043
rect 311216 3012 312093 3040
rect 311216 3000 311222 3012
rect 312081 3009 312093 3012
rect 312127 3009 312139 3043
rect 312081 3003 312139 3009
rect 314838 3000 314844 3052
rect 314896 3040 314902 3052
rect 315942 3040 315948 3052
rect 314896 3012 315948 3040
rect 314896 3000 314902 3012
rect 315942 3000 315948 3012
rect 316000 3000 316006 3052
rect 317966 3000 317972 3052
rect 318024 3040 318030 3052
rect 333514 3040 333520 3052
rect 318024 3012 333520 3040
rect 318024 3000 318030 3012
rect 333514 3000 333520 3012
rect 333572 3000 333578 3052
rect 356790 3000 356796 3052
rect 356848 3040 356854 3052
rect 417878 3040 417884 3052
rect 356848 3012 417884 3040
rect 356848 3000 356854 3012
rect 417878 3000 417884 3012
rect 417936 3000 417942 3052
rect 311084 2944 312768 2972
rect 260374 2864 260380 2916
rect 260432 2904 260438 2916
rect 312630 2904 312636 2916
rect 260432 2876 312636 2904
rect 260432 2864 260438 2876
rect 312630 2864 312636 2876
rect 312688 2864 312694 2916
rect 284662 2796 284668 2848
rect 284720 2836 284726 2848
rect 312078 2836 312084 2848
rect 284720 2808 312084 2836
rect 284720 2796 284726 2808
rect 312078 2796 312084 2808
rect 312136 2796 312142 2848
rect 312740 2836 312768 2944
rect 315574 2932 315580 2984
rect 315632 2972 315638 2984
rect 375558 2972 375564 2984
rect 315632 2944 375564 2972
rect 315632 2932 315638 2944
rect 375558 2932 375564 2944
rect 375616 2932 375622 2984
rect 314286 2864 314292 2916
rect 314344 2904 314350 2916
rect 354214 2904 354220 2916
rect 314344 2876 354220 2904
rect 314344 2864 314350 2876
rect 354214 2864 354220 2876
rect 354272 2864 354278 2916
rect 364242 2864 364248 2916
rect 364300 2904 364306 2916
rect 421006 2904 421012 2916
rect 364300 2876 421012 2904
rect 364300 2864 364306 2876
rect 421006 2864 421012 2876
rect 421064 2864 421070 2916
rect 315758 2836 315764 2848
rect 312740 2808 315764 2836
rect 315758 2796 315764 2808
rect 315816 2796 315822 2848
rect 357342 2796 357348 2848
rect 357400 2836 357406 2848
rect 390646 2836 390652 2848
rect 357400 2808 390652 2836
rect 357400 2796 357406 2808
rect 390646 2796 390652 2808
rect 390704 2796 390710 2848
<< via1 >>
rect 369860 617516 369912 617568
rect 371148 617516 371200 617568
rect 463700 617516 463752 617568
rect 464988 617516 465040 617568
rect 494060 617516 494112 617568
rect 495348 617516 495400 617568
rect 3424 616836 3476 616888
rect 134524 616836 134576 616888
rect 22836 616768 22888 616820
rect 23388 616768 23440 616820
rect 34980 616768 35032 616820
rect 35808 616768 35860 616820
rect 53012 616768 53064 616820
rect 53748 616768 53800 616820
rect 77300 616768 77352 616820
rect 78496 616768 78548 616820
rect 113732 616768 113784 616820
rect 114376 616768 114428 616820
rect 143908 616768 143960 616820
rect 299204 616768 299256 616820
rect 310612 616768 310664 616820
rect 311808 616768 311860 616820
rect 313372 616768 313424 616820
rect 428740 616768 428792 616820
rect 4620 616700 4672 616752
rect 5448 616700 5500 616752
rect 65156 616700 65208 616752
rect 66168 616700 66220 616752
rect 80428 616700 80480 616752
rect 81348 616700 81400 616752
rect 114100 616700 114152 616752
rect 265164 616700 265216 616752
rect 285312 616700 285364 616752
rect 462044 616700 462096 616752
rect 471060 616700 471112 616752
rect 471888 616700 471940 616752
rect 106740 616632 106792 616684
rect 125876 616632 125928 616684
rect 131764 616632 131816 616684
rect 315396 616632 315448 616684
rect 392308 616632 392360 616684
rect 393228 616632 393280 616684
rect 101588 616564 101640 616616
rect 322204 616564 322256 616616
rect 356060 616564 356112 616616
rect 382556 616564 382608 616616
rect 36360 616496 36412 616548
rect 134892 616496 134944 616548
rect 137836 616496 137888 616548
rect 363604 616496 363656 616548
rect 17224 616428 17276 616480
rect 128820 616428 128872 616480
rect 153844 616428 153896 616480
rect 183284 616428 183336 616480
rect 184572 616428 184624 616480
rect 416596 616428 416648 616480
rect 71228 616360 71280 616412
rect 314108 616360 314160 616412
rect 331772 616360 331824 616412
rect 371792 616360 371844 616412
rect 389824 616360 389876 616412
rect 443828 616360 443880 616412
rect 110604 616292 110656 616344
rect 425704 616292 425756 616344
rect 6828 616224 6880 616276
rect 122748 616224 122800 616276
rect 136548 616224 136600 616276
rect 452844 616224 452896 616276
rect 9864 616156 9916 616208
rect 25780 616156 25832 616208
rect 28908 616156 28960 616208
rect 103520 616156 103572 616208
rect 104532 616156 104584 616208
rect 438308 616156 438360 616208
rect 1676 616088 1728 616140
rect 359464 616088 359516 616140
rect 395344 616088 395396 616140
rect 468116 616088 468168 616140
rect 78588 616020 78640 616072
rect 162124 616020 162176 616072
rect 222660 616020 222712 616072
rect 83372 615952 83424 616004
rect 160744 615952 160796 616004
rect 233424 616020 233476 616072
rect 277308 616020 277360 616072
rect 281356 616020 281408 616072
rect 404452 616020 404504 616072
rect 314016 615952 314068 616004
rect 95516 615884 95568 615936
rect 167736 615884 167788 615936
rect 262036 615884 262088 615936
rect 346492 615884 346544 615936
rect 98460 615816 98512 615868
rect 153200 615816 153252 615868
rect 216220 615816 216272 615868
rect 289268 615816 289320 615868
rect 143816 615748 143868 615800
rect 198556 615748 198608 615800
rect 210516 615748 210568 615800
rect 211068 615748 211120 615800
rect 247592 615748 247644 615800
rect 298468 615748 298520 615800
rect 268384 615680 268436 615732
rect 313556 615680 313608 615732
rect 280252 615544 280304 615596
rect 281448 615544 281500 615596
rect 334716 615544 334768 615596
rect 492956 615476 493008 615528
rect 364248 614975 364300 614984
rect 364248 614941 364257 614975
rect 364257 614941 364291 614975
rect 364291 614941 364300 614975
rect 364248 614932 364300 614941
rect 137192 613844 137244 613896
rect 167276 613887 167328 613896
rect 167276 613853 167285 613887
rect 167285 613853 167319 613887
rect 167319 613853 167328 613887
rect 167276 613844 167328 613853
rect 175740 613912 175792 613964
rect 167644 613887 167696 613896
rect 167644 613853 167653 613887
rect 167653 613853 167687 613887
rect 167687 613853 167696 613887
rect 167644 613844 167696 613853
rect 175648 613776 175700 613828
rect 167920 613751 167972 613760
rect 167920 613717 167929 613751
rect 167929 613717 167963 613751
rect 167963 613717 167972 613751
rect 167920 613708 167972 613717
rect 182088 612756 182140 612808
rect 495440 612756 495492 612808
rect 402428 611668 402480 611720
rect 237840 611532 237892 611584
rect 283012 610623 283064 610632
rect 283012 610589 283021 610623
rect 283021 610589 283055 610623
rect 283055 610589 283064 610623
rect 283012 610580 283064 610589
rect 435272 610580 435324 610632
rect 283288 610555 283340 610564
rect 283288 610521 283297 610555
rect 283297 610521 283331 610555
rect 283331 610521 283340 610555
rect 283288 610512 283340 610521
rect 283380 610555 283432 610564
rect 283380 610521 283389 610555
rect 283389 610521 283423 610555
rect 283423 610521 283432 610555
rect 283380 610512 283432 610521
rect 456800 610512 456852 610564
rect 440884 610444 440936 610496
rect 434904 610240 434956 610292
rect 283012 610172 283064 610224
rect 419540 610172 419592 610224
rect 386420 609492 386472 609544
rect 480260 608812 480312 608864
rect 3056 608744 3108 608796
rect 6184 608744 6236 608796
rect 334900 607971 334952 607980
rect 334900 607937 334909 607971
rect 334909 607937 334943 607971
rect 334943 607937 334952 607971
rect 334900 607928 334952 607937
rect 334716 607767 334768 607776
rect 334716 607733 334725 607767
rect 334725 607733 334759 607767
rect 334759 607733 334768 607767
rect 334716 607724 334768 607733
rect 236460 607316 236512 607368
rect 263876 607180 263928 607232
rect 228456 606883 228508 606892
rect 228456 606849 228490 606883
rect 228490 606849 228508 606883
rect 228456 606840 228508 606849
rect 310796 606636 310848 606688
rect 231860 606432 231912 606484
rect 3424 604460 3476 604512
rect 55496 604460 55548 604512
rect 78496 604052 78548 604104
rect 184572 601443 184624 601452
rect 184572 601409 184581 601443
rect 184581 601409 184615 601443
rect 184615 601409 184624 601443
rect 184572 601400 184624 601409
rect 196440 600788 196492 600840
rect 23020 600763 23072 600772
rect 23020 600729 23054 600763
rect 23054 600729 23072 600763
rect 23020 600720 23072 600729
rect 142436 600652 142488 600704
rect 233424 600287 233476 600296
rect 233424 600253 233433 600287
rect 233433 600253 233467 600287
rect 233467 600253 233476 600287
rect 233424 600244 233476 600253
rect 3516 599292 3568 599344
rect 53840 599360 53892 599412
rect 50160 599063 50212 599072
rect 50160 599029 50169 599063
rect 50169 599029 50203 599063
rect 50203 599029 50212 599063
rect 50160 599020 50212 599029
rect 331220 599224 331272 599276
rect 158904 599156 158956 599208
rect 158996 599088 159048 599140
rect 79232 599020 79284 599072
rect 325608 599020 325660 599072
rect 314200 598952 314252 599004
rect 495440 598952 495492 599004
rect 247592 596683 247644 596692
rect 247592 596649 247601 596683
rect 247601 596649 247635 596683
rect 247635 596649 247644 596683
rect 247592 596640 247644 596649
rect 206008 596547 206060 596556
rect 206008 596513 206017 596547
rect 206017 596513 206051 596547
rect 206051 596513 206060 596547
rect 206008 596504 206060 596513
rect 205456 596343 205508 596352
rect 205456 596309 205465 596343
rect 205465 596309 205499 596343
rect 205499 596309 205508 596343
rect 205456 596300 205508 596309
rect 205824 596343 205876 596352
rect 205824 596309 205833 596343
rect 205833 596309 205867 596343
rect 205867 596309 205876 596343
rect 205824 596300 205876 596309
rect 205916 596343 205968 596352
rect 205916 596309 205925 596343
rect 205925 596309 205959 596343
rect 205959 596309 205968 596343
rect 205916 596300 205968 596309
rect 2780 595008 2832 595060
rect 5172 595008 5224 595060
rect 492956 591243 493008 591252
rect 492956 591209 492965 591243
rect 492965 591209 492999 591243
rect 492999 591209 493008 591243
rect 492956 591200 493008 591209
rect 494336 591039 494388 591048
rect 494336 591005 494345 591039
rect 494345 591005 494379 591039
rect 494379 591005 494388 591039
rect 494336 590996 494388 591005
rect 111892 590928 111944 590980
rect 419540 590631 419592 590640
rect 419540 590597 419549 590631
rect 419549 590597 419583 590631
rect 419583 590597 419592 590631
rect 419540 590588 419592 590597
rect 419356 590563 419408 590572
rect 419356 590529 419365 590563
rect 419365 590529 419399 590563
rect 419399 590529 419408 590563
rect 419356 590520 419408 590529
rect 435364 590520 435416 590572
rect 419632 590359 419684 590368
rect 419632 590325 419641 590359
rect 419641 590325 419675 590359
rect 419675 590325 419684 590359
rect 419632 590316 419684 590325
rect 463424 587299 463476 587308
rect 463424 587265 463433 587299
rect 463433 587265 463467 587299
rect 463467 587265 463476 587299
rect 463424 587256 463476 587265
rect 463516 587299 463568 587308
rect 463516 587265 463525 587299
rect 463525 587265 463559 587299
rect 463559 587265 463568 587299
rect 463516 587256 463568 587265
rect 495532 587256 495584 587308
rect 463148 587231 463200 587240
rect 463148 587197 463157 587231
rect 463157 587197 463191 587231
rect 463191 587197 463200 587231
rect 463148 587188 463200 587197
rect 203984 587052 204036 587104
rect 416688 586848 416740 586900
rect 2780 586508 2832 586560
rect 4896 586508 4948 586560
rect 313372 586211 313424 586220
rect 313372 586177 313381 586211
rect 313381 586177 313415 586211
rect 313415 586177 313424 586211
rect 313372 586168 313424 586177
rect 4804 585556 4856 585608
rect 106740 584715 106792 584724
rect 106740 584681 106749 584715
rect 106749 584681 106783 584715
rect 106783 584681 106792 584715
rect 106740 584672 106792 584681
rect 206008 584400 206060 584452
rect 262496 584400 262548 584452
rect 142068 583992 142120 584044
rect 201500 583967 201552 583976
rect 201500 583933 201509 583967
rect 201509 583933 201543 583967
rect 201543 583933 201552 583967
rect 201500 583924 201552 583933
rect 206008 583856 206060 583908
rect 201960 583831 202012 583840
rect 201960 583797 201969 583831
rect 201969 583797 202003 583831
rect 202003 583797 202012 583831
rect 201960 583788 202012 583797
rect 405924 583423 405976 583432
rect 405924 583389 405933 583423
rect 405933 583389 405967 583423
rect 405967 583389 405976 583423
rect 405924 583380 405976 583389
rect 28908 580728 28960 580780
rect 482652 580703 482704 580712
rect 482652 580669 482661 580703
rect 482661 580669 482695 580703
rect 482695 580669 482704 580703
rect 482652 580660 482704 580669
rect 482744 580703 482796 580712
rect 482744 580669 482753 580703
rect 482753 580669 482787 580703
rect 482787 580669 482796 580703
rect 482744 580660 482796 580669
rect 372712 580524 372764 580576
rect 291200 579028 291252 579080
rect 121368 578892 121420 578944
rect 180432 578688 180484 578740
rect 396724 578935 396776 578944
rect 396724 578901 396733 578935
rect 396733 578901 396767 578935
rect 396767 578901 396776 578935
rect 396724 578892 396776 578901
rect 403440 578892 403492 578944
rect 482744 578892 482796 578944
rect 3608 578348 3660 578400
rect 2780 577260 2832 577312
rect 4988 577260 5040 577312
rect 247684 576920 247736 576972
rect 233332 576852 233384 576904
rect 423588 576895 423640 576904
rect 423588 576861 423597 576895
rect 423597 576861 423631 576895
rect 423631 576861 423640 576895
rect 423588 576852 423640 576861
rect 66168 576172 66220 576224
rect 43076 572704 43128 572756
rect 495440 572704 495492 572756
rect 231860 572092 231912 572144
rect 196440 572067 196492 572076
rect 196440 572033 196449 572067
rect 196449 572033 196483 572067
rect 196483 572033 196492 572067
rect 196440 572024 196492 572033
rect 422944 572024 422996 572076
rect 213828 571888 213880 571940
rect 445668 571820 445720 571872
rect 236460 571115 236512 571124
rect 236460 571081 236469 571115
rect 236469 571081 236503 571115
rect 236503 571081 236512 571115
rect 236460 571072 236512 571081
rect 237564 570979 237616 570988
rect 237564 570945 237582 570979
rect 237582 570945 237616 570979
rect 237564 570936 237616 570945
rect 237840 570979 237892 570988
rect 237840 570945 237849 570979
rect 237849 570945 237883 570979
rect 237883 570945 237892 570979
rect 237840 570936 237892 570945
rect 285312 570979 285364 570988
rect 285312 570945 285321 570979
rect 285321 570945 285355 570979
rect 285355 570945 285364 570979
rect 285312 570936 285364 570945
rect 236460 570732 236512 570784
rect 417884 570732 417936 570784
rect 376484 569279 376536 569288
rect 376484 569245 376493 569279
rect 376493 569245 376527 569279
rect 376527 569245 376536 569279
rect 376484 569236 376536 569245
rect 473728 567103 473780 567112
rect 473728 567069 473737 567103
rect 473737 567069 473771 567103
rect 473771 567069 473780 567103
rect 473728 567060 473780 567069
rect 473912 567103 473964 567112
rect 473912 567069 473921 567103
rect 473921 567069 473955 567103
rect 473955 567069 473964 567103
rect 473912 567060 473964 567069
rect 451924 566924 451976 566976
rect 78588 566219 78640 566228
rect 78588 566185 78597 566219
rect 78597 566185 78631 566219
rect 78631 566185 78640 566219
rect 78588 566176 78640 566185
rect 233700 565972 233752 566024
rect 325608 566015 325660 566024
rect 325608 565981 325617 566015
rect 325617 565981 325651 566015
rect 325651 565981 325660 566015
rect 325608 565972 325660 565981
rect 325792 566015 325844 566024
rect 325792 565981 325801 566015
rect 325801 565981 325835 566015
rect 325835 565981 325844 566015
rect 325792 565972 325844 565981
rect 75920 565904 75972 565956
rect 76288 565947 76340 565956
rect 76288 565913 76297 565947
rect 76297 565913 76331 565947
rect 76331 565913 76340 565947
rect 76288 565904 76340 565913
rect 208308 565904 208360 565956
rect 325516 565947 325568 565956
rect 325516 565913 325525 565947
rect 325525 565913 325559 565947
rect 325559 565913 325568 565947
rect 325516 565904 325568 565913
rect 158444 565836 158496 565888
rect 15016 561731 15068 561740
rect 15016 561697 15025 561731
rect 15025 561697 15059 561731
rect 15059 561697 15068 561731
rect 15016 561688 15068 561697
rect 51448 561688 51500 561740
rect 15292 561663 15344 561672
rect 15292 561629 15301 561663
rect 15301 561629 15335 561663
rect 15335 561629 15344 561663
rect 15292 561620 15344 561629
rect 258908 561620 258960 561672
rect 123392 561552 123444 561604
rect 203984 559147 204036 559156
rect 203984 559113 203993 559147
rect 203993 559113 204027 559147
rect 204027 559113 204036 559147
rect 203984 559104 204036 559113
rect 255688 558968 255740 559020
rect 2872 558900 2924 558952
rect 101404 558900 101456 558952
rect 204352 558943 204404 558952
rect 204352 558909 204361 558943
rect 204361 558909 204395 558943
rect 204395 558909 204404 558943
rect 204352 558900 204404 558909
rect 403440 557379 403492 557388
rect 403440 557345 403449 557379
rect 403449 557345 403483 557379
rect 403483 557345 403492 557379
rect 403440 557336 403492 557345
rect 82728 557132 82780 557184
rect 327264 556928 327316 556980
rect 403348 557175 403400 557184
rect 403348 557141 403357 557175
rect 403357 557141 403391 557175
rect 403391 557141 403400 557175
rect 403348 557132 403400 557141
rect 331496 556792 331548 556844
rect 310612 556724 310664 556776
rect 316684 556656 316736 556708
rect 403440 556180 403492 556232
rect 406016 556180 406068 556232
rect 313924 555092 313976 555144
rect 2780 554752 2832 554804
rect 6276 554752 6328 554804
rect 316776 554752 316828 554804
rect 495440 554752 495492 554804
rect 330852 554047 330904 554056
rect 330852 554013 330861 554047
rect 330861 554013 330895 554047
rect 330895 554013 330904 554047
rect 330852 554004 330904 554013
rect 268292 553528 268344 553580
rect 268568 553571 268620 553580
rect 268568 553537 268577 553571
rect 268577 553537 268611 553571
rect 268611 553537 268620 553571
rect 268752 553571 268804 553580
rect 268568 553528 268620 553537
rect 268752 553537 268760 553571
rect 268760 553537 268794 553571
rect 268794 553537 268804 553571
rect 268752 553528 268804 553537
rect 268844 553571 268896 553580
rect 268844 553537 268853 553571
rect 268853 553537 268887 553571
rect 268887 553537 268896 553571
rect 268844 553528 268896 553537
rect 447784 553460 447836 553512
rect 376208 553392 376260 553444
rect 434904 551871 434956 551880
rect 434904 551837 434908 551871
rect 434908 551837 434942 551871
rect 434942 551837 434956 551871
rect 434904 551828 434956 551837
rect 435272 551871 435324 551880
rect 435272 551837 435280 551871
rect 435280 551837 435314 551871
rect 435314 551837 435324 551871
rect 435272 551828 435324 551837
rect 435364 551871 435416 551880
rect 435364 551837 435373 551871
rect 435373 551837 435407 551871
rect 435407 551837 435416 551871
rect 435364 551828 435416 551837
rect 434996 551803 435048 551812
rect 434996 551769 435005 551803
rect 435005 551769 435039 551803
rect 435039 551769 435048 551803
rect 434996 551760 435048 551769
rect 435088 551803 435140 551812
rect 435088 551769 435097 551803
rect 435097 551769 435131 551803
rect 435131 551769 435140 551803
rect 435088 551760 435140 551769
rect 434720 551735 434772 551744
rect 434720 551701 434729 551735
rect 434729 551701 434763 551735
rect 434763 551701 434772 551735
rect 434720 551692 434772 551701
rect 311164 549244 311216 549296
rect 495440 549244 495492 549296
rect 231860 548675 231912 548684
rect 231860 548641 231869 548675
rect 231869 548641 231903 548675
rect 231903 548641 231912 548675
rect 231860 548632 231912 548641
rect 260656 548564 260708 548616
rect 232136 548539 232188 548548
rect 232136 548505 232170 548539
rect 232170 548505 232188 548539
rect 232136 548496 232188 548505
rect 279240 548496 279292 548548
rect 343640 548496 343692 548548
rect 380624 547519 380676 547528
rect 380624 547485 380633 547519
rect 380633 547485 380667 547519
rect 380667 547485 380676 547519
rect 380624 547476 380676 547485
rect 119528 547408 119580 547460
rect 379244 547383 379296 547392
rect 379244 547349 379253 547383
rect 379253 547349 379287 547383
rect 379287 547349 379296 547383
rect 379244 547340 379296 547349
rect 121828 546839 121880 546848
rect 121828 546805 121837 546839
rect 121837 546805 121871 546839
rect 121871 546805 121880 546839
rect 121828 546796 121880 546805
rect 3148 545096 3200 545148
rect 265072 545096 265124 545148
rect 363512 545096 363564 545148
rect 495440 545096 495492 545148
rect 3424 544212 3476 544264
rect 416596 544255 416648 544264
rect 416596 544221 416605 544255
rect 416605 544221 416639 544255
rect 416639 544221 416648 544255
rect 416596 544212 416648 544221
rect 334716 543804 334768 543856
rect 157248 543779 157300 543788
rect 157248 543745 157257 543779
rect 157257 543745 157291 543779
rect 157291 543745 157300 543779
rect 157248 543736 157300 543745
rect 157432 543779 157484 543788
rect 157432 543745 157441 543779
rect 157441 543745 157475 543779
rect 157475 543745 157484 543779
rect 157432 543736 157484 543745
rect 157524 543736 157576 543788
rect 469588 543736 469640 543788
rect 330852 542308 330904 542360
rect 495440 542308 495492 542360
rect 119528 541739 119580 541748
rect 119528 541705 119537 541739
rect 119537 541705 119571 541739
rect 119571 541705 119580 541739
rect 119528 541696 119580 541705
rect 123300 541628 123352 541680
rect 120080 541535 120132 541544
rect 120080 541501 120089 541535
rect 120089 541501 120123 541535
rect 120123 541501 120132 541535
rect 120080 541492 120132 541501
rect 379244 541560 379296 541612
rect 367744 541492 367796 541544
rect 119988 541467 120040 541476
rect 119988 541433 119997 541467
rect 119997 541433 120031 541467
rect 120031 541433 120040 541467
rect 119988 541424 120040 541433
rect 2872 540948 2924 541000
rect 388444 540948 388496 541000
rect 158444 540515 158496 540524
rect 158444 540481 158453 540515
rect 158453 540481 158487 540515
rect 158487 540481 158496 540515
rect 158444 540472 158496 540481
rect 158628 540515 158680 540524
rect 158628 540481 158637 540515
rect 158637 540481 158671 540515
rect 158671 540481 158680 540515
rect 158628 540472 158680 540481
rect 221464 540404 221516 540456
rect 158720 540336 158772 540388
rect 158812 540336 158864 540388
rect 159088 540379 159140 540388
rect 159088 540345 159097 540379
rect 159097 540345 159131 540379
rect 159131 540345 159140 540379
rect 159088 540336 159140 540345
rect 158628 540268 158680 540320
rect 273904 540268 273956 540320
rect 462320 539520 462372 539572
rect 463148 539520 463200 539572
rect 59452 539427 59504 539436
rect 59452 539393 59461 539427
rect 59461 539393 59495 539427
rect 59495 539393 59504 539427
rect 59452 539384 59504 539393
rect 463424 539384 463476 539436
rect 462320 539316 462372 539368
rect 326344 539248 326396 539300
rect 59176 539223 59228 539232
rect 59176 539189 59185 539223
rect 59185 539189 59219 539223
rect 59219 539189 59228 539223
rect 59176 539180 59228 539189
rect 59636 539223 59688 539232
rect 59636 539189 59645 539223
rect 59645 539189 59679 539223
rect 59679 539189 59688 539223
rect 59636 539180 59688 539189
rect 6368 537684 6420 537736
rect 229008 537684 229060 537736
rect 3148 536800 3200 536852
rect 6736 536800 6788 536852
rect 176936 536800 176988 536852
rect 495440 536800 495492 536852
rect 3516 536596 3568 536648
rect 404268 534692 404320 534744
rect 473912 534692 473964 534744
rect 331496 534667 331548 534676
rect 331496 534633 331505 534667
rect 331505 534633 331539 534667
rect 331539 534633 331548 534667
rect 331496 534624 331548 534633
rect 331312 534463 331364 534472
rect 331312 534429 331321 534463
rect 331321 534429 331355 534463
rect 331355 534429 331364 534463
rect 331312 534420 331364 534429
rect 334900 534420 334952 534472
rect 331496 534284 331548 534336
rect 402980 534284 403032 534336
rect 404268 534284 404320 534336
rect 361488 533944 361540 533996
rect 4528 533740 4580 533792
rect 430764 533740 430816 533792
rect 342444 531607 342496 531616
rect 342444 531573 342453 531607
rect 342453 531573 342487 531607
rect 342487 531573 342496 531607
rect 342444 531564 342496 531573
rect 355600 529023 355652 529032
rect 355600 528989 355609 529023
rect 355609 528989 355643 529023
rect 355643 528989 355652 529023
rect 355600 528980 355652 528989
rect 417976 528980 418028 529032
rect 355508 528887 355560 528896
rect 355508 528853 355517 528887
rect 355517 528853 355551 528887
rect 355551 528853 355560 528887
rect 355508 528844 355560 528853
rect 121828 528504 121880 528556
rect 495440 528504 495492 528556
rect 81348 528300 81400 528352
rect 12992 527935 13044 527944
rect 12992 527901 13001 527935
rect 13001 527901 13035 527935
rect 13035 527901 13044 527935
rect 12992 527892 13044 527901
rect 353944 527935 353996 527944
rect 353944 527901 353953 527935
rect 353953 527901 353987 527935
rect 353987 527901 353996 527935
rect 353944 527892 353996 527901
rect 12716 527867 12768 527876
rect 12716 527833 12734 527867
rect 12734 527833 12768 527867
rect 12716 527824 12768 527833
rect 417792 527756 417844 527808
rect 112536 527416 112588 527468
rect 380624 527416 380676 527468
rect 375656 527255 375708 527264
rect 375656 527221 375665 527255
rect 375665 527221 375699 527255
rect 375699 527221 375708 527255
rect 375656 527212 375708 527221
rect 380624 527144 380676 527196
rect 383660 527144 383712 527196
rect 273628 526328 273680 526380
rect 121000 526167 121052 526176
rect 121000 526133 121009 526167
rect 121009 526133 121043 526167
rect 121043 526133 121052 526167
rect 121000 526124 121052 526133
rect 158720 526124 158772 526176
rect 262772 525283 262824 525292
rect 262772 525249 262781 525283
rect 262781 525249 262815 525283
rect 262815 525249 262824 525283
rect 262772 525240 262824 525249
rect 262496 525215 262548 525224
rect 262496 525181 262505 525215
rect 262505 525181 262539 525215
rect 262539 525181 262548 525215
rect 262496 525172 262548 525181
rect 262680 525215 262732 525224
rect 262680 525181 262689 525215
rect 262689 525181 262723 525215
rect 262723 525181 262732 525215
rect 262680 525172 262732 525181
rect 290832 525172 290884 525224
rect 351460 525215 351512 525224
rect 351460 525181 351469 525215
rect 351469 525181 351503 525215
rect 351503 525181 351512 525215
rect 351460 525172 351512 525181
rect 351736 525215 351788 525224
rect 351736 525181 351745 525215
rect 351745 525181 351779 525215
rect 351779 525181 351788 525215
rect 351736 525172 351788 525181
rect 452108 525172 452160 525224
rect 15292 525036 15344 525088
rect 153476 525036 153528 525088
rect 158628 524764 158680 524816
rect 75920 524696 75972 524748
rect 351736 524739 351788 524748
rect 351736 524705 351745 524739
rect 351745 524705 351779 524739
rect 351779 524705 351788 524739
rect 351736 524696 351788 524705
rect 27436 524560 27488 524612
rect 157524 524560 157576 524612
rect 11428 524535 11480 524544
rect 11428 524501 11437 524535
rect 11437 524501 11471 524535
rect 11471 524501 11480 524535
rect 11428 524492 11480 524501
rect 113088 524492 113140 524544
rect 291108 518755 291160 518764
rect 291108 518721 291117 518755
rect 291117 518721 291151 518755
rect 291151 518721 291160 518755
rect 291108 518712 291160 518721
rect 289820 518644 289872 518696
rect 290832 518576 290884 518628
rect 244924 518508 244976 518560
rect 319904 514879 319956 514888
rect 319904 514845 319913 514879
rect 319913 514845 319947 514879
rect 319947 514845 319956 514879
rect 319904 514836 319956 514845
rect 435088 514836 435140 514888
rect 3332 514768 3384 514820
rect 14464 514768 14516 514820
rect 319812 514811 319864 514820
rect 319812 514777 319821 514811
rect 319821 514777 319855 514811
rect 319855 514777 319864 514811
rect 319812 514768 319864 514777
rect 309692 514360 309744 514412
rect 267648 514292 267700 514344
rect 405832 514335 405884 514344
rect 405832 514301 405841 514335
rect 405841 514301 405875 514335
rect 405875 514301 405884 514335
rect 405832 514292 405884 514301
rect 406016 514335 406068 514344
rect 406016 514301 406025 514335
rect 406025 514301 406059 514335
rect 406059 514301 406068 514335
rect 406016 514292 406068 514301
rect 409604 514292 409656 514344
rect 157248 514156 157300 514208
rect 405372 514199 405424 514208
rect 405372 514165 405381 514199
rect 405381 514165 405415 514199
rect 405415 514165 405424 514199
rect 405372 514156 405424 514165
rect 328460 513952 328512 514004
rect 7840 513680 7892 513732
rect 46020 513791 46072 513800
rect 46020 513757 46029 513791
rect 46029 513757 46063 513791
rect 46063 513757 46072 513791
rect 260656 513859 260708 513868
rect 260656 513825 260665 513859
rect 260665 513825 260699 513859
rect 260699 513825 260708 513859
rect 260656 513816 260708 513825
rect 276940 513816 276992 513868
rect 46020 513748 46072 513757
rect 46204 513723 46256 513732
rect 46204 513689 46213 513723
rect 46213 513689 46247 513723
rect 46247 513689 46256 513723
rect 46204 513680 46256 513689
rect 177028 513680 177080 513732
rect 410524 513748 410576 513800
rect 45744 513655 45796 513664
rect 45744 513621 45753 513655
rect 45753 513621 45787 513655
rect 45787 513621 45796 513655
rect 45744 513612 45796 513621
rect 259184 513612 259236 513664
rect 317328 510935 317380 510944
rect 317328 510901 317337 510935
rect 317337 510901 317371 510935
rect 317371 510901 317380 510935
rect 317328 510892 317380 510901
rect 8024 509260 8076 509312
rect 495440 509260 495492 509312
rect 326344 508011 326396 508020
rect 326344 507977 326353 508011
rect 326353 507977 326387 508011
rect 326387 507977 326396 508011
rect 326344 507968 326396 507977
rect 496360 507900 496412 507952
rect 59176 507832 59228 507884
rect 426624 507875 426676 507884
rect 426624 507841 426633 507875
rect 426633 507841 426667 507875
rect 426667 507841 426676 507875
rect 426624 507832 426676 507841
rect 426808 507875 426860 507884
rect 426808 507841 426817 507875
rect 426817 507841 426851 507875
rect 426851 507841 426860 507875
rect 426808 507832 426860 507841
rect 324964 507807 325016 507816
rect 324964 507773 324973 507807
rect 324973 507773 325007 507807
rect 325007 507773 325016 507807
rect 324964 507764 325016 507773
rect 324964 507628 325016 507680
rect 383936 507628 383988 507680
rect 426900 507671 426952 507680
rect 426900 507637 426909 507671
rect 426909 507637 426943 507671
rect 426943 507637 426952 507671
rect 426900 507628 426952 507637
rect 247684 507467 247736 507476
rect 247684 507433 247693 507467
rect 247693 507433 247727 507467
rect 247727 507433 247736 507467
rect 247684 507424 247736 507433
rect 247592 507263 247644 507272
rect 247592 507229 247601 507263
rect 247601 507229 247635 507263
rect 247635 507229 247644 507263
rect 247592 507220 247644 507229
rect 41788 507152 41840 507204
rect 496360 507220 496412 507272
rect 373816 507152 373868 507204
rect 248144 507127 248196 507136
rect 248144 507093 248153 507127
rect 248153 507093 248187 507127
rect 248187 507093 248196 507127
rect 248144 507084 248196 507093
rect 3148 505112 3200 505164
rect 349804 505112 349856 505164
rect 384028 504568 384080 504620
rect 406568 504568 406620 504620
rect 383844 504407 383896 504416
rect 383844 504373 383853 504407
rect 383853 504373 383887 504407
rect 383887 504373 383896 504407
rect 383844 504364 383896 504373
rect 443092 504364 443144 504416
rect 406568 503684 406620 503736
rect 464160 503684 464212 503736
rect 153844 502188 153896 502240
rect 421012 500828 421064 500880
rect 420736 500803 420788 500812
rect 420736 500769 420745 500803
rect 420745 500769 420779 500803
rect 420779 500769 420788 500803
rect 420736 500760 420788 500769
rect 420920 500735 420972 500744
rect 420920 500701 420929 500735
rect 420929 500701 420963 500735
rect 420963 500701 420972 500735
rect 420920 500692 420972 500701
rect 420552 500667 420604 500676
rect 420552 500633 420561 500667
rect 420561 500633 420595 500667
rect 420595 500633 420604 500667
rect 420552 500624 420604 500633
rect 420644 500667 420696 500676
rect 420644 500633 420653 500667
rect 420653 500633 420687 500667
rect 420687 500633 420696 500667
rect 420644 500624 420696 500633
rect 369124 500556 369176 500608
rect 481824 500624 481876 500676
rect 190368 500055 190420 500064
rect 190368 500021 190377 500055
rect 190377 500021 190411 500055
rect 190411 500021 190420 500055
rect 190368 500012 190420 500021
rect 208308 498108 208360 498160
rect 208584 498083 208636 498092
rect 208584 498049 208593 498083
rect 208593 498049 208627 498083
rect 208627 498049 208636 498083
rect 208584 498040 208636 498049
rect 233792 498040 233844 498092
rect 208308 497836 208360 497888
rect 331588 497836 331640 497888
rect 2780 496952 2832 497004
rect 5356 496952 5408 497004
rect 255596 496383 255648 496392
rect 255596 496349 255605 496383
rect 255605 496349 255639 496383
rect 255639 496349 255648 496383
rect 255596 496340 255648 496349
rect 351460 496204 351512 496256
rect 255688 495907 255740 495916
rect 255688 495873 255697 495907
rect 255697 495873 255731 495907
rect 255731 495873 255740 495907
rect 255688 495864 255740 495873
rect 255596 495796 255648 495848
rect 380716 495864 380768 495916
rect 423588 496068 423640 496120
rect 290280 495796 290332 495848
rect 6460 494572 6512 494624
rect 3700 494164 3752 494216
rect 29644 493144 29696 493196
rect 93768 493144 93820 493196
rect 32312 493051 32364 493060
rect 32312 493017 32321 493051
rect 32321 493017 32355 493051
rect 32355 493017 32364 493051
rect 32312 493008 32364 493017
rect 32404 492983 32456 492992
rect 32404 492949 32413 492983
rect 32413 492949 32447 492983
rect 32447 492949 32456 492983
rect 32772 492983 32824 492992
rect 32404 492940 32456 492949
rect 32772 492949 32781 492983
rect 32781 492949 32815 492983
rect 32815 492949 32824 492983
rect 32772 492940 32824 492949
rect 276940 492192 276992 492244
rect 276940 492099 276992 492108
rect 276940 492065 276949 492099
rect 276949 492065 276983 492099
rect 276983 492065 276992 492099
rect 276940 492056 276992 492065
rect 208492 492031 208544 492040
rect 208492 491997 208501 492031
rect 208501 491997 208535 492031
rect 208535 491997 208544 492031
rect 208492 491988 208544 491997
rect 237380 491988 237432 492040
rect 277308 491920 277360 491972
rect 324964 491988 325016 492040
rect 207112 491895 207164 491904
rect 207112 491861 207121 491895
rect 207121 491861 207155 491895
rect 207155 491861 207164 491895
rect 384304 491920 384356 491972
rect 207112 491852 207164 491861
rect 429292 491852 429344 491904
rect 277308 491648 277360 491700
rect 378784 491648 378836 491700
rect 367008 491580 367060 491632
rect 237380 489812 237432 489864
rect 238208 489812 238260 489864
rect 276940 489812 276992 489864
rect 412916 489855 412968 489864
rect 412916 489821 412925 489855
rect 412925 489821 412959 489855
rect 412959 489821 412968 489855
rect 412916 489812 412968 489821
rect 432512 489812 432564 489864
rect 248328 489787 248380 489796
rect 248328 489753 248362 489787
rect 248362 489753 248380 489787
rect 248328 489744 248380 489753
rect 249432 489719 249484 489728
rect 249432 489685 249441 489719
rect 249441 489685 249475 489719
rect 249475 489685 249484 489719
rect 249432 489676 249484 489685
rect 27528 489472 27580 489524
rect 414296 489719 414348 489728
rect 414296 489685 414305 489719
rect 414305 489685 414339 489719
rect 414339 489685 414348 489719
rect 414296 489676 414348 489685
rect 423956 489676 424008 489728
rect 470048 489175 470100 489184
rect 470048 489141 470057 489175
rect 470057 489141 470091 489175
rect 470091 489141 470100 489175
rect 470048 489132 470100 489141
rect 21640 487296 21692 487348
rect 9588 487228 9640 487280
rect 237656 487228 237708 487280
rect 417792 487228 417844 487280
rect 417884 487228 417936 487280
rect 7104 487160 7156 487212
rect 417976 487203 418028 487212
rect 417976 487169 417985 487203
rect 417985 487169 418019 487203
rect 418019 487169 418028 487203
rect 417976 487160 418028 487169
rect 422024 487160 422076 487212
rect 29644 487024 29696 487076
rect 264060 485639 264112 485648
rect 264060 485605 264069 485639
rect 264069 485605 264103 485639
rect 264103 485605 264112 485639
rect 264060 485596 264112 485605
rect 263692 485528 263744 485580
rect 420736 485528 420788 485580
rect 263876 485503 263928 485512
rect 263876 485469 263885 485503
rect 263885 485469 263919 485503
rect 263919 485469 263928 485503
rect 263876 485460 263928 485469
rect 420552 485460 420604 485512
rect 263508 485367 263560 485376
rect 263508 485333 263517 485367
rect 263517 485333 263551 485367
rect 263551 485333 263560 485367
rect 263508 485324 263560 485333
rect 263692 485367 263744 485376
rect 263692 485333 263701 485367
rect 263701 485333 263735 485367
rect 263735 485333 263744 485367
rect 263692 485324 263744 485333
rect 263784 485367 263836 485376
rect 263784 485333 263793 485367
rect 263793 485333 263827 485367
rect 263827 485333 263836 485367
rect 264152 485392 264204 485444
rect 477776 485392 477828 485444
rect 263784 485324 263836 485333
rect 421012 485324 421064 485376
rect 464160 484075 464212 484084
rect 464160 484041 464169 484075
rect 464169 484041 464203 484075
rect 464203 484041 464212 484075
rect 464160 484032 464212 484041
rect 464252 484075 464304 484084
rect 464252 484041 464261 484075
rect 464261 484041 464295 484075
rect 464295 484041 464304 484075
rect 464252 484032 464304 484041
rect 463976 483939 464028 483948
rect 463976 483905 463985 483939
rect 463985 483905 464019 483939
rect 464019 483905 464028 483939
rect 463976 483896 464028 483905
rect 464344 483939 464396 483948
rect 464344 483905 464353 483939
rect 464353 483905 464387 483939
rect 464387 483905 464396 483939
rect 464344 483896 464396 483905
rect 167276 483760 167328 483812
rect 382556 482443 382608 482452
rect 382556 482409 382565 482443
rect 382565 482409 382599 482443
rect 382599 482409 382608 482443
rect 382556 482400 382608 482409
rect 383936 482307 383988 482316
rect 383936 482273 383945 482307
rect 383945 482273 383979 482307
rect 383979 482273 383988 482307
rect 383936 482264 383988 482273
rect 412916 482196 412968 482248
rect 383752 482060 383804 482112
rect 22836 480632 22888 480684
rect 327724 480564 327776 480616
rect 16212 480471 16264 480480
rect 16212 480437 16221 480471
rect 16221 480437 16255 480471
rect 16255 480437 16264 480471
rect 16212 480428 16264 480437
rect 238208 480131 238260 480140
rect 238208 480097 238217 480131
rect 238217 480097 238251 480131
rect 238251 480097 238260 480131
rect 238208 480088 238260 480097
rect 238484 479995 238536 480004
rect 238484 479961 238518 479995
rect 238518 479961 238536 479995
rect 238484 479952 238536 479961
rect 259368 479884 259420 479936
rect 2780 479000 2832 479052
rect 5264 479000 5316 479052
rect 259368 478864 259420 478916
rect 331680 478864 331732 478916
rect 360568 475736 360620 475788
rect 297640 475668 297692 475720
rect 495532 475711 495584 475720
rect 495532 475677 495541 475711
rect 495541 475677 495575 475711
rect 495575 475677 495584 475711
rect 495532 475668 495584 475677
rect 495624 475711 495676 475720
rect 495624 475677 495633 475711
rect 495633 475677 495667 475711
rect 495667 475677 495676 475711
rect 495624 475668 495676 475677
rect 5908 475532 5960 475584
rect 9772 475328 9824 475380
rect 194600 475328 194652 475380
rect 93768 473628 93820 473680
rect 112444 473560 112496 473612
rect 93768 473492 93820 473544
rect 97080 473492 97132 473544
rect 228916 473492 228968 473544
rect 93308 473356 93360 473408
rect 93676 473356 93728 473408
rect 203064 473399 203116 473408
rect 203064 473365 203073 473399
rect 203073 473365 203107 473399
rect 203107 473365 203116 473399
rect 203064 473356 203116 473365
rect 263508 471316 263560 471368
rect 198280 471291 198332 471300
rect 198280 471257 198289 471291
rect 198289 471257 198323 471291
rect 198323 471257 198332 471291
rect 198280 471248 198332 471257
rect 198464 471291 198516 471300
rect 198464 471257 198473 471291
rect 198473 471257 198507 471291
rect 198507 471257 198516 471291
rect 198464 471248 198516 471257
rect 268844 471248 268896 471300
rect 194784 470908 194836 470960
rect 344284 470840 344336 470892
rect 384028 470636 384080 470688
rect 432512 469820 432564 469872
rect 443920 469820 443972 469872
rect 494336 469820 494388 469872
rect 167920 469752 167972 469804
rect 8944 469548 8996 469600
rect 463976 469548 464028 469600
rect 315764 469208 315816 469260
rect 495440 469208 495492 469260
rect 334624 467440 334676 467492
rect 112996 467372 113048 467424
rect 247592 467372 247644 467424
rect 111892 467211 111944 467220
rect 111892 467177 111901 467211
rect 111901 467177 111935 467211
rect 111935 467177 111944 467211
rect 111892 467168 111944 467177
rect 194784 467168 194836 467220
rect 208492 467168 208544 467220
rect 112996 467032 113048 467084
rect 112628 466964 112680 467016
rect 112812 466896 112864 466948
rect 195060 466939 195112 466948
rect 195060 466905 195094 466939
rect 195094 466905 195112 466939
rect 195060 466896 195112 466905
rect 340880 466828 340932 466880
rect 207204 465400 207256 465452
rect 224408 465375 224460 465384
rect 120080 465196 120132 465248
rect 224408 465341 224417 465375
rect 224417 465341 224451 465375
rect 224451 465341 224460 465375
rect 224408 465332 224460 465341
rect 255596 465264 255648 465316
rect 311900 465196 311952 465248
rect 338028 463700 338080 463752
rect 6552 463020 6604 463072
rect 3332 460912 3384 460964
rect 170404 460955 170456 460964
rect 170404 460921 170413 460955
rect 170413 460921 170447 460955
rect 170447 460921 170456 460955
rect 170404 460912 170456 460921
rect 358084 460912 358136 460964
rect 356704 457580 356756 457632
rect 254216 457215 254268 457224
rect 254216 457181 254225 457215
rect 254225 457181 254259 457215
rect 254259 457181 254268 457215
rect 254216 457172 254268 457181
rect 254124 457079 254176 457088
rect 254124 457045 254133 457079
rect 254133 457045 254167 457079
rect 254167 457045 254176 457079
rect 254124 457036 254176 457045
rect 484216 455404 484268 455456
rect 495440 455404 495492 455456
rect 314292 454316 314344 454368
rect 315304 453271 315356 453280
rect 315304 453237 315313 453271
rect 315313 453237 315347 453271
rect 315347 453237 315356 453271
rect 315304 453228 315356 453237
rect 43168 451256 43220 451308
rect 333520 451324 333572 451376
rect 54024 451299 54076 451308
rect 54024 451265 54033 451299
rect 54033 451265 54067 451299
rect 54067 451265 54076 451299
rect 54024 451256 54076 451265
rect 53472 451095 53524 451104
rect 53472 451061 53481 451095
rect 53481 451061 53515 451095
rect 53515 451061 53524 451095
rect 53472 451052 53524 451061
rect 53932 451095 53984 451104
rect 53932 451061 53941 451095
rect 53941 451061 53975 451095
rect 53975 451061 53984 451095
rect 53932 451052 53984 451061
rect 142344 448536 142396 448588
rect 175740 448468 175792 448520
rect 176016 448511 176068 448520
rect 176016 448477 176025 448511
rect 176025 448477 176059 448511
rect 176059 448477 176068 448511
rect 176016 448468 176068 448477
rect 419356 448468 419408 448520
rect 175556 448443 175608 448452
rect 175556 448409 175565 448443
rect 175565 448409 175599 448443
rect 175599 448409 175608 448443
rect 175556 448400 175608 448409
rect 175648 448443 175700 448452
rect 175648 448409 175657 448443
rect 175657 448409 175691 448443
rect 175691 448409 175700 448443
rect 175648 448400 175700 448409
rect 178316 448400 178368 448452
rect 383844 448332 383896 448384
rect 64788 447831 64840 447840
rect 64788 447797 64797 447831
rect 64797 447797 64831 447831
rect 64831 447797 64840 447831
rect 64788 447788 64840 447797
rect 53472 446904 53524 446956
rect 112260 446947 112312 446956
rect 112260 446913 112269 446947
rect 112269 446913 112303 446947
rect 112303 446913 112312 446947
rect 112260 446904 112312 446913
rect 112352 446947 112404 446956
rect 112352 446913 112361 446947
rect 112361 446913 112395 446947
rect 112395 446913 112404 446947
rect 112352 446904 112404 446913
rect 112444 446879 112496 446888
rect 112444 446845 112453 446879
rect 112453 446845 112487 446879
rect 112487 446845 112496 446879
rect 112444 446836 112496 446845
rect 140780 446836 140832 446888
rect 383936 446836 383988 446888
rect 88340 446700 88392 446752
rect 333520 446743 333572 446752
rect 333520 446709 333529 446743
rect 333529 446709 333563 446743
rect 333563 446709 333572 446743
rect 333520 446700 333572 446709
rect 152372 443683 152424 443692
rect 152372 443649 152381 443683
rect 152381 443649 152415 443683
rect 152415 443649 152424 443683
rect 152372 443640 152424 443649
rect 423864 443640 423916 443692
rect 152464 443615 152516 443624
rect 152464 443581 152473 443615
rect 152473 443581 152507 443615
rect 152507 443581 152516 443615
rect 152464 443572 152516 443581
rect 224408 443572 224460 443624
rect 112628 443436 112680 443488
rect 424048 443479 424100 443488
rect 424048 443445 424057 443479
rect 424057 443445 424091 443479
rect 424091 443445 424100 443479
rect 424048 443436 424100 443445
rect 152280 443096 152332 443148
rect 153016 443003 153068 443012
rect 153016 442969 153025 443003
rect 153025 442969 153059 443003
rect 153059 442969 153068 443003
rect 153016 442960 153068 442969
rect 281356 442595 281408 442604
rect 281356 442561 281365 442595
rect 281365 442561 281399 442595
rect 281399 442561 281408 442595
rect 281356 442552 281408 442561
rect 376208 441983 376260 441992
rect 376208 441949 376217 441983
rect 376217 441949 376251 441983
rect 376251 441949 376260 441983
rect 376208 441940 376260 441949
rect 376116 441847 376168 441856
rect 376116 441813 376125 441847
rect 376125 441813 376159 441847
rect 376159 441813 376168 441847
rect 376116 441804 376168 441813
rect 311348 441600 311400 441652
rect 495440 441600 495492 441652
rect 412088 439832 412140 439884
rect 336556 439764 336608 439816
rect 195244 439696 195296 439748
rect 412272 439696 412324 439748
rect 418804 439807 418856 439816
rect 418804 439773 418813 439807
rect 418813 439773 418847 439807
rect 418847 439773 418856 439807
rect 418804 439764 418856 439773
rect 418988 439671 419040 439680
rect 418988 439637 418997 439671
rect 418997 439637 419031 439671
rect 419031 439637 419040 439671
rect 418988 439628 419040 439637
rect 43168 439424 43220 439476
rect 41788 439331 41840 439340
rect 41788 439297 41797 439331
rect 41797 439297 41831 439331
rect 41831 439297 41840 439331
rect 41788 439288 41840 439297
rect 281448 436908 281500 436960
rect 420644 435072 420696 435124
rect 47676 435004 47728 435056
rect 44088 434868 44140 434920
rect 48044 434979 48096 434988
rect 48044 434945 48053 434979
rect 48053 434945 48087 434979
rect 48087 434945 48096 434979
rect 48044 434936 48096 434945
rect 48228 434979 48280 434988
rect 48228 434945 48237 434979
rect 48237 434945 48271 434979
rect 48271 434945 48280 434979
rect 48228 434936 48280 434945
rect 48136 434868 48188 434920
rect 143080 434868 143132 434920
rect 47860 434843 47912 434852
rect 47860 434809 47869 434843
rect 47869 434809 47903 434843
rect 47903 434809 47912 434843
rect 47860 434800 47912 434809
rect 263692 434800 263744 434852
rect 436744 434732 436796 434784
rect 91468 434299 91520 434308
rect 91468 434265 91477 434299
rect 91477 434265 91511 434299
rect 91511 434265 91520 434299
rect 91468 434256 91520 434265
rect 293684 434256 293736 434308
rect 159088 434188 159140 434240
rect 267740 433372 267792 433424
rect 3332 433304 3384 433356
rect 338764 433304 338816 433356
rect 281356 432191 281408 432200
rect 281356 432157 281365 432191
rect 281365 432157 281399 432191
rect 281399 432157 281408 432191
rect 281356 432148 281408 432157
rect 308312 432148 308364 432200
rect 281632 432123 281684 432132
rect 281632 432089 281666 432123
rect 281666 432089 281684 432123
rect 281632 432080 281684 432089
rect 282736 432055 282788 432064
rect 282736 432021 282745 432055
rect 282745 432021 282779 432055
rect 282779 432021 282788 432055
rect 282736 432012 282788 432021
rect 496544 432012 496596 432064
rect 133696 429496 133748 429548
rect 142436 429539 142488 429548
rect 142436 429505 142445 429539
rect 142445 429505 142479 429539
rect 142479 429505 142488 429539
rect 142436 429496 142488 429505
rect 142344 429403 142396 429412
rect 142344 429369 142353 429403
rect 142353 429369 142387 429403
rect 142387 429369 142396 429403
rect 142344 429360 142396 429369
rect 412272 428451 412324 428460
rect 412272 428417 412281 428451
rect 412281 428417 412315 428451
rect 412315 428417 412324 428451
rect 412272 428408 412324 428417
rect 412364 428451 412416 428460
rect 412364 428417 412373 428451
rect 412373 428417 412407 428451
rect 412407 428417 412416 428451
rect 412364 428408 412416 428417
rect 290004 428340 290056 428392
rect 184572 428204 184624 428256
rect 412088 428247 412140 428256
rect 412088 428213 412097 428247
rect 412097 428213 412131 428247
rect 412131 428213 412140 428247
rect 412088 428204 412140 428213
rect 311808 426708 311860 426760
rect 3332 425144 3384 425196
rect 6644 425144 6696 425196
rect 91468 425076 91520 425128
rect 92388 425076 92440 425128
rect 95884 425076 95936 425128
rect 239036 424532 239088 424584
rect 46020 424464 46072 424516
rect 449900 424532 449952 424584
rect 312084 424464 312136 424516
rect 312084 423648 312136 423700
rect 495992 423648 496044 423700
rect 15016 423512 15068 423564
rect 331404 423555 331456 423564
rect 132592 423444 132644 423496
rect 133696 423487 133748 423496
rect 133696 423453 133705 423487
rect 133705 423453 133739 423487
rect 133739 423453 133748 423487
rect 133696 423444 133748 423453
rect 133880 423487 133932 423496
rect 133880 423453 133888 423487
rect 133888 423453 133922 423487
rect 133922 423453 133932 423487
rect 133880 423444 133932 423453
rect 133972 423487 134024 423496
rect 133972 423453 133981 423487
rect 133981 423453 134015 423487
rect 134015 423453 134024 423487
rect 133972 423444 134024 423453
rect 134156 423444 134208 423496
rect 331404 423521 331413 423555
rect 331413 423521 331447 423555
rect 331447 423521 331456 423555
rect 331404 423512 331456 423521
rect 331220 423444 331272 423496
rect 331496 423487 331548 423496
rect 331496 423453 331505 423487
rect 331505 423453 331539 423487
rect 331539 423453 331548 423487
rect 331496 423444 331548 423453
rect 331680 423487 331732 423496
rect 331680 423453 331689 423487
rect 331689 423453 331723 423487
rect 331723 423453 331732 423487
rect 331680 423444 331732 423453
rect 89260 423308 89312 423360
rect 134340 423351 134392 423360
rect 134340 423317 134349 423351
rect 134349 423317 134383 423351
rect 134383 423317 134392 423351
rect 134340 423308 134392 423317
rect 244464 423376 244516 423428
rect 385132 423376 385184 423428
rect 27528 423147 27580 423156
rect 27528 423113 27537 423147
rect 27537 423113 27571 423147
rect 27571 423113 27580 423147
rect 27528 423104 27580 423113
rect 133972 423104 134024 423156
rect 205272 423104 205324 423156
rect 451464 423104 451516 423156
rect 134156 423036 134208 423088
rect 205364 423036 205416 423088
rect 27436 423011 27488 423020
rect 27436 422977 27445 423011
rect 27445 422977 27479 423011
rect 27479 422977 27488 423011
rect 27436 422968 27488 422977
rect 92388 422968 92440 423020
rect 121000 422900 121052 422952
rect 67364 422832 67416 422884
rect 55404 422764 55456 422816
rect 9680 422560 9732 422612
rect 133880 422560 133932 422612
rect 443920 421311 443972 421320
rect 443920 421277 443929 421311
rect 443929 421277 443963 421311
rect 443963 421277 443972 421311
rect 443920 421268 443972 421277
rect 470416 421268 470468 421320
rect 338212 421200 338264 421252
rect 442540 421175 442592 421184
rect 442540 421141 442549 421175
rect 442549 421141 442583 421175
rect 442583 421141 442592 421175
rect 442540 421132 442592 421141
rect 3976 417528 4028 417580
rect 334072 417571 334124 417580
rect 334072 417537 334081 417571
rect 334081 417537 334115 417571
rect 334115 417537 334124 417571
rect 334072 417528 334124 417537
rect 334348 417503 334400 417512
rect 334348 417469 334357 417503
rect 334357 417469 334391 417503
rect 334391 417469 334400 417503
rect 334348 417460 334400 417469
rect 203064 417392 203116 417444
rect 5080 417324 5132 417376
rect 136548 417163 136600 417172
rect 136548 417129 136557 417163
rect 136557 417129 136591 417163
rect 136591 417129 136600 417163
rect 136548 417120 136600 417129
rect 152464 415488 152516 415540
rect 101496 415420 101548 415472
rect 279240 415395 279292 415404
rect 279240 415361 279249 415395
rect 279249 415361 279283 415395
rect 279283 415361 279292 415395
rect 279240 415352 279292 415361
rect 8116 415284 8168 415336
rect 257068 415327 257120 415336
rect 257068 415293 257077 415327
rect 257077 415293 257111 415327
rect 257111 415293 257120 415327
rect 257068 415284 257120 415293
rect 262496 415284 262548 415336
rect 232136 415216 232188 415268
rect 279608 415327 279660 415336
rect 279608 415293 279617 415327
rect 279617 415293 279651 415327
rect 279651 415293 279660 415327
rect 346860 415420 346912 415472
rect 346584 415352 346636 415404
rect 279608 415284 279660 415293
rect 95608 415148 95660 415200
rect 119620 414783 119672 414792
rect 119620 414749 119629 414783
rect 119629 414749 119663 414783
rect 119663 414749 119672 414783
rect 119620 414740 119672 414749
rect 318064 414264 318116 414316
rect 402428 414239 402480 414248
rect 402428 414205 402437 414239
rect 402437 414205 402471 414239
rect 402471 414205 402480 414239
rect 402428 414196 402480 414205
rect 403808 414103 403860 414112
rect 403808 414069 403817 414103
rect 403817 414069 403851 414103
rect 403851 414069 403860 414103
rect 403808 414060 403860 414069
rect 485596 414060 485648 414112
rect 258908 413899 258960 413908
rect 258908 413865 258917 413899
rect 258917 413865 258951 413899
rect 258951 413865 258960 413899
rect 258908 413856 258960 413865
rect 281356 413652 281408 413704
rect 205640 413584 205692 413636
rect 143816 412811 143868 412820
rect 143816 412777 143825 412811
rect 143825 412777 143859 412811
rect 143859 412777 143868 412811
rect 143816 412768 143868 412777
rect 254124 412632 254176 412684
rect 257436 412632 257488 412684
rect 389180 411884 389232 411936
rect 4068 411476 4120 411528
rect 99656 411043 99708 411052
rect 99656 411009 99665 411043
rect 99665 411009 99699 411043
rect 99699 411009 99708 411043
rect 99656 411000 99708 411009
rect 99840 411043 99892 411052
rect 99840 411009 99849 411043
rect 99849 411009 99883 411043
rect 99883 411009 99892 411043
rect 99840 411000 99892 411009
rect 254124 410932 254176 410984
rect 112536 410635 112588 410644
rect 112536 410601 112545 410635
rect 112545 410601 112579 410635
rect 112579 410601 112588 410635
rect 112536 410592 112588 410601
rect 112996 410635 113048 410644
rect 112996 410601 113005 410635
rect 113005 410601 113039 410635
rect 113039 410601 113048 410635
rect 112996 410592 113048 410601
rect 325792 410864 325844 410916
rect 335544 410592 335596 410644
rect 99840 410524 99892 410576
rect 331496 410524 331548 410576
rect 113088 410499 113140 410508
rect 113088 410465 113097 410499
rect 113097 410465 113131 410499
rect 113131 410465 113140 410499
rect 113088 410456 113140 410465
rect 112812 410431 112864 410440
rect 112812 410397 112821 410431
rect 112821 410397 112855 410431
rect 112855 410397 112864 410431
rect 112812 410388 112864 410397
rect 375380 410388 375432 410440
rect 375656 410388 375708 410440
rect 112812 410252 112864 410304
rect 253112 410320 253164 410372
rect 55312 409955 55364 409964
rect 55312 409921 55321 409955
rect 55321 409921 55355 409955
rect 55355 409921 55364 409955
rect 55312 409912 55364 409921
rect 55496 409955 55548 409964
rect 55496 409921 55505 409955
rect 55505 409921 55539 409955
rect 55539 409921 55548 409955
rect 55496 409912 55548 409921
rect 198464 409912 198516 409964
rect 89444 409844 89496 409896
rect 57152 409411 57204 409420
rect 57152 409377 57161 409411
rect 57161 409377 57195 409411
rect 57195 409377 57204 409411
rect 57152 409368 57204 409377
rect 57336 409368 57388 409420
rect 342904 409368 342956 409420
rect 56876 409343 56928 409352
rect 56876 409309 56885 409343
rect 56885 409309 56919 409343
rect 56919 409309 56928 409343
rect 56876 409300 56928 409309
rect 56692 409207 56744 409216
rect 56692 409173 56701 409207
rect 56701 409173 56735 409207
rect 56735 409173 56744 409207
rect 56692 409164 56744 409173
rect 177304 409300 177356 409352
rect 92296 409232 92348 409284
rect 56876 408960 56928 409012
rect 90640 409164 90692 409216
rect 3332 407124 3384 407176
rect 11704 407124 11756 407176
rect 316868 407124 316920 407176
rect 495440 407124 495492 407176
rect 3332 406988 3384 407040
rect 4068 406988 4120 407040
rect 35808 406036 35860 406088
rect 114100 405603 114152 405612
rect 114100 405569 114109 405603
rect 114109 405569 114143 405603
rect 114143 405569 114152 405603
rect 114100 405560 114152 405569
rect 3056 403180 3108 403232
rect 170404 402908 170456 402960
rect 495440 402908 495492 402960
rect 119988 401684 120040 401736
rect 2964 401616 3016 401668
rect 312176 401616 312228 401668
rect 414296 400664 414348 400716
rect 67088 400639 67140 400648
rect 67088 400605 67097 400639
rect 67097 400605 67131 400639
rect 67131 400605 67140 400639
rect 67088 400596 67140 400605
rect 67364 400639 67416 400648
rect 67364 400605 67373 400639
rect 67373 400605 67407 400639
rect 67407 400605 67416 400639
rect 67364 400596 67416 400605
rect 67456 400639 67508 400648
rect 67456 400605 67465 400639
rect 67465 400605 67499 400639
rect 67499 400605 67508 400639
rect 67456 400596 67508 400605
rect 67640 400596 67692 400648
rect 423772 400596 423824 400648
rect 283288 400528 283340 400580
rect 67640 400503 67692 400512
rect 67640 400469 67649 400503
rect 67649 400469 67683 400503
rect 67683 400469 67692 400503
rect 67640 400460 67692 400469
rect 314384 399916 314436 399968
rect 375472 399508 375524 399560
rect 376116 399508 376168 399560
rect 253112 399415 253164 399424
rect 253112 399381 253121 399415
rect 253121 399381 253155 399415
rect 253155 399381 253164 399415
rect 253112 399372 253164 399381
rect 426716 399372 426768 399424
rect 400036 398463 400088 398472
rect 400036 398429 400045 398463
rect 400045 398429 400079 398463
rect 400079 398429 400088 398463
rect 400036 398420 400088 398429
rect 326528 397783 326580 397792
rect 326528 397749 326537 397783
rect 326537 397749 326571 397783
rect 326571 397749 326580 397783
rect 326528 397740 326580 397749
rect 316960 397536 317012 397588
rect 495440 397536 495492 397588
rect 211068 397468 211120 397520
rect 398104 396244 398156 396296
rect 43076 395811 43128 395820
rect 43076 395777 43085 395811
rect 43085 395777 43119 395811
rect 43119 395777 43128 395811
rect 43076 395768 43128 395777
rect 3792 395564 3844 395616
rect 380624 395224 380676 395276
rect 11796 395199 11848 395208
rect 11796 395165 11805 395199
rect 11805 395165 11839 395199
rect 11839 395165 11848 395199
rect 11796 395156 11848 395165
rect 380716 395199 380768 395208
rect 380716 395165 380725 395199
rect 380725 395165 380759 395199
rect 380759 395165 380768 395199
rect 380716 395156 380768 395165
rect 380900 395063 380952 395072
rect 380900 395029 380909 395063
rect 380909 395029 380943 395063
rect 380943 395029 380952 395063
rect 380900 395020 380952 395029
rect 433984 395020 434036 395072
rect 22836 394859 22888 394868
rect 22836 394825 22845 394859
rect 22845 394825 22879 394859
rect 22879 394825 22888 394859
rect 22836 394816 22888 394825
rect 22928 394680 22980 394732
rect 45744 394748 45796 394800
rect 360384 394680 360436 394732
rect 452108 394179 452160 394188
rect 452108 394145 452117 394179
rect 452117 394145 452151 394179
rect 452151 394145 452160 394179
rect 452108 394136 452160 394145
rect 451924 394111 451976 394120
rect 451924 394077 451933 394111
rect 451933 394077 451967 394111
rect 451967 394077 451976 394111
rect 451924 394068 451976 394077
rect 167828 393728 167880 393780
rect 451556 393975 451608 393984
rect 451556 393941 451565 393975
rect 451565 393941 451599 393975
rect 451599 393941 451608 393975
rect 451556 393932 451608 393941
rect 6092 393388 6144 393440
rect 330484 392300 330536 392352
rect 3608 389648 3660 389700
rect 3792 389648 3844 389700
rect 3608 389172 3660 389224
rect 214564 389172 214616 389224
rect 346768 387651 346820 387660
rect 346768 387617 346777 387651
rect 346777 387617 346811 387651
rect 346811 387617 346820 387651
rect 346768 387608 346820 387617
rect 346860 387651 346912 387660
rect 346860 387617 346869 387651
rect 346869 387617 346903 387651
rect 346903 387617 346912 387651
rect 346860 387608 346912 387617
rect 346492 387583 346544 387592
rect 346492 387549 346501 387583
rect 346501 387549 346535 387583
rect 346535 387549 346544 387583
rect 346492 387540 346544 387549
rect 346584 387583 346636 387592
rect 346584 387549 346593 387583
rect 346593 387549 346627 387583
rect 346627 387549 346636 387583
rect 346584 387540 346636 387549
rect 450452 387540 450504 387592
rect 407396 387472 407448 387524
rect 346308 387447 346360 387456
rect 346308 387413 346317 387447
rect 346317 387413 346351 387447
rect 346351 387413 346360 387447
rect 346308 387404 346360 387413
rect 367744 387107 367796 387116
rect 367744 387073 367753 387107
rect 367753 387073 367787 387107
rect 367787 387073 367796 387107
rect 367744 387064 367796 387073
rect 371240 387064 371292 387116
rect 22100 386996 22152 387048
rect 368388 386996 368440 387048
rect 412272 387132 412324 387184
rect 367560 386971 367612 386980
rect 367560 386937 367569 386971
rect 367569 386937 367603 386971
rect 367603 386937 367612 386971
rect 367560 386928 367612 386937
rect 368020 386903 368072 386912
rect 368020 386869 368029 386903
rect 368029 386869 368063 386903
rect 368063 386869 368072 386903
rect 368020 386860 368072 386869
rect 450636 386860 450688 386912
rect 353944 384956 353996 385008
rect 495440 384956 495492 385008
rect 95976 384752 96028 384804
rect 108304 384727 108356 384736
rect 108304 384693 108313 384727
rect 108313 384693 108347 384727
rect 108347 384693 108356 384727
rect 108304 384684 108356 384693
rect 89444 384523 89496 384532
rect 89444 384489 89453 384523
rect 89453 384489 89487 384523
rect 89487 384489 89496 384523
rect 89444 384480 89496 384489
rect 414388 384412 414440 384464
rect 89260 384387 89312 384396
rect 89260 384353 89269 384387
rect 89269 384353 89303 384387
rect 89303 384353 89312 384387
rect 89260 384344 89312 384353
rect 142436 384344 142488 384396
rect 132592 384319 132644 384328
rect 88800 384251 88852 384260
rect 88800 384217 88809 384251
rect 88809 384217 88843 384251
rect 88843 384217 88852 384251
rect 88800 384208 88852 384217
rect 132592 384285 132601 384319
rect 132601 384285 132635 384319
rect 132635 384285 132644 384319
rect 132592 384276 132644 384285
rect 403808 384276 403860 384328
rect 200488 384208 200540 384260
rect 232688 384208 232740 384260
rect 89076 384183 89128 384192
rect 89076 384149 89085 384183
rect 89085 384149 89119 384183
rect 89119 384149 89128 384183
rect 89076 384140 89128 384149
rect 89168 384183 89220 384192
rect 89168 384149 89177 384183
rect 89177 384149 89211 384183
rect 89211 384149 89220 384183
rect 89168 384140 89220 384149
rect 103520 384183 103572 384192
rect 103520 384149 103529 384183
rect 103529 384149 103563 384183
rect 103563 384149 103572 384183
rect 132408 384183 132460 384192
rect 103520 384140 103572 384149
rect 132408 384149 132417 384183
rect 132417 384149 132451 384183
rect 132451 384149 132460 384183
rect 132408 384140 132460 384149
rect 177028 383979 177080 383988
rect 177028 383945 177037 383979
rect 177037 383945 177071 383979
rect 177071 383945 177080 383979
rect 177028 383936 177080 383945
rect 259184 383936 259236 383988
rect 177212 383843 177264 383852
rect 177212 383809 177221 383843
rect 177221 383809 177255 383843
rect 177255 383809 177264 383843
rect 177212 383800 177264 383809
rect 177304 383843 177356 383852
rect 177304 383809 177313 383843
rect 177313 383809 177347 383843
rect 177347 383809 177356 383843
rect 177304 383800 177356 383809
rect 199660 383800 199712 383852
rect 199752 383732 199804 383784
rect 279608 383868 279660 383920
rect 200120 383775 200172 383784
rect 200120 383741 200129 383775
rect 200129 383741 200163 383775
rect 200163 383741 200172 383775
rect 334072 383800 334124 383852
rect 200120 383732 200172 383741
rect 311992 383732 312044 383784
rect 317052 383664 317104 383716
rect 199660 383596 199712 383648
rect 13728 383188 13780 383240
rect 130384 383231 130436 383240
rect 130384 383197 130393 383231
rect 130393 383197 130427 383231
rect 130427 383197 130436 383231
rect 130384 383188 130436 383197
rect 322296 383231 322348 383240
rect 322296 383197 322305 383231
rect 322305 383197 322339 383231
rect 322339 383197 322348 383231
rect 322296 383188 322348 383197
rect 136548 381488 136600 381540
rect 464344 381488 464396 381540
rect 39396 381012 39448 381064
rect 39396 380919 39448 380928
rect 39396 380885 39405 380919
rect 39405 380885 39439 380919
rect 39439 380885 39448 380919
rect 39396 380876 39448 380885
rect 40592 380876 40644 380928
rect 89260 381012 89312 381064
rect 136088 380876 136140 380928
rect 136548 380876 136600 380928
rect 274456 380443 274508 380452
rect 274456 380409 274465 380443
rect 274465 380409 274499 380443
rect 274499 380409 274508 380443
rect 274456 380400 274508 380409
rect 71872 378879 71924 378888
rect 71872 378845 71881 378879
rect 71881 378845 71915 378879
rect 71915 378845 71924 378879
rect 71872 378836 71924 378845
rect 259552 378836 259604 378888
rect 95792 378768 95844 378820
rect 70584 378743 70636 378752
rect 70584 378709 70593 378743
rect 70593 378709 70627 378743
rect 70627 378709 70636 378743
rect 70584 378700 70636 378709
rect 309692 375819 309744 375828
rect 309692 375785 309701 375819
rect 309701 375785 309735 375819
rect 309735 375785 309744 375819
rect 309692 375776 309744 375785
rect 308312 375683 308364 375692
rect 308312 375649 308321 375683
rect 308321 375649 308355 375683
rect 308355 375649 308364 375683
rect 308312 375640 308364 375649
rect 5356 375572 5408 375624
rect 342260 375572 342312 375624
rect 8852 375504 8904 375556
rect 309692 375436 309744 375488
rect 366732 375436 366784 375488
rect 409420 375139 409472 375148
rect 409420 375105 409429 375139
rect 409429 375105 409463 375139
rect 409463 375105 409472 375139
rect 409420 375096 409472 375105
rect 405004 375028 405056 375080
rect 409604 375071 409656 375080
rect 409604 375037 409613 375071
rect 409613 375037 409647 375071
rect 409647 375037 409656 375071
rect 409604 375028 409656 375037
rect 419080 375028 419132 375080
rect 409052 374935 409104 374944
rect 409052 374901 409061 374935
rect 409061 374901 409095 374935
rect 409095 374901 409104 374935
rect 409052 374892 409104 374901
rect 95608 374731 95660 374740
rect 95608 374697 95617 374731
rect 95617 374697 95651 374731
rect 95651 374697 95660 374731
rect 95608 374688 95660 374697
rect 450452 374731 450504 374740
rect 450452 374697 450461 374731
rect 450461 374697 450495 374731
rect 450495 374697 450504 374731
rect 450452 374688 450504 374697
rect 95976 374595 96028 374604
rect 95976 374561 95985 374595
rect 95985 374561 96019 374595
rect 96019 374561 96028 374595
rect 95976 374552 96028 374561
rect 95792 374527 95844 374536
rect 95792 374493 95801 374527
rect 95801 374493 95835 374527
rect 95835 374493 95844 374527
rect 95792 374484 95844 374493
rect 152372 374484 152424 374536
rect 450636 374527 450688 374536
rect 450636 374493 450645 374527
rect 450645 374493 450679 374527
rect 450679 374493 450688 374527
rect 450636 374484 450688 374493
rect 441988 372351 442040 372360
rect 441988 372317 441997 372351
rect 441997 372317 442031 372351
rect 442031 372317 442040 372351
rect 441988 372308 442040 372317
rect 233700 371875 233752 371884
rect 233700 371841 233709 371875
rect 233709 371841 233743 371875
rect 233743 371841 233752 371875
rect 233700 371832 233752 371841
rect 233792 371671 233844 371680
rect 233792 371637 233801 371671
rect 233801 371637 233835 371671
rect 233835 371637 233844 371671
rect 233792 371628 233844 371637
rect 366824 371628 366876 371680
rect 214748 370175 214800 370184
rect 214748 370141 214757 370175
rect 214757 370141 214791 370175
rect 214791 370141 214800 370175
rect 214748 370132 214800 370141
rect 293684 369087 293736 369096
rect 293684 369053 293693 369087
rect 293693 369053 293727 369087
rect 293727 369053 293736 369087
rect 293684 369044 293736 369053
rect 325516 369044 325568 369096
rect 335636 369112 335688 369164
rect 311624 368908 311676 368960
rect 2780 366664 2832 366716
rect 4712 366664 4764 366716
rect 360568 366571 360620 366580
rect 360568 366537 360577 366571
rect 360577 366537 360611 366571
rect 360611 366537 360620 366571
rect 360568 366528 360620 366537
rect 360384 366435 360436 366444
rect 360384 366401 360393 366435
rect 360393 366401 360427 366435
rect 360427 366401 360436 366435
rect 360384 366392 360436 366401
rect 360200 366367 360252 366376
rect 360200 366333 360209 366367
rect 360209 366333 360243 366367
rect 360243 366333 360252 366367
rect 360200 366324 360252 366333
rect 314568 365712 314620 365764
rect 495440 365712 495492 365764
rect 473728 365483 473780 365492
rect 143080 365372 143132 365424
rect 473728 365449 473737 365483
rect 473737 365449 473771 365483
rect 473771 365449 473780 365483
rect 473728 365440 473780 365449
rect 263876 365372 263928 365424
rect 264060 365304 264112 365356
rect 473636 365347 473688 365356
rect 473636 365313 473645 365347
rect 473645 365313 473679 365347
rect 473679 365313 473688 365347
rect 473636 365304 473688 365313
rect 143080 365100 143132 365152
rect 355600 365100 355652 365152
rect 470416 364735 470468 364744
rect 470416 364701 470425 364735
rect 470425 364701 470459 364735
rect 470459 364701 470468 364735
rect 470416 364692 470468 364701
rect 486976 364692 487028 364744
rect 248144 364624 248196 364676
rect 496360 364556 496412 364608
rect 153016 362584 153068 362636
rect 180432 362627 180484 362636
rect 180432 362593 180441 362627
rect 180441 362593 180475 362627
rect 180475 362593 180484 362627
rect 180432 362584 180484 362593
rect 180064 362491 180116 362500
rect 180064 362457 180073 362491
rect 180073 362457 180107 362491
rect 180107 362457 180116 362491
rect 180064 362448 180116 362457
rect 316040 362516 316092 362568
rect 426992 361564 427044 361616
rect 495440 361564 495492 361616
rect 244372 360383 244424 360392
rect 244372 360349 244381 360383
rect 244381 360349 244415 360383
rect 244415 360349 244424 360383
rect 244372 360340 244424 360349
rect 402796 360383 402848 360392
rect 402796 360349 402805 360383
rect 402805 360349 402839 360383
rect 402839 360349 402848 360383
rect 402796 360340 402848 360349
rect 402980 360383 403032 360392
rect 402980 360349 402989 360383
rect 402989 360349 403023 360383
rect 403023 360349 403032 360383
rect 402980 360340 403032 360349
rect 336188 360204 336240 360256
rect 361488 359907 361540 359916
rect 361488 359873 361497 359907
rect 361497 359873 361531 359907
rect 361531 359873 361540 359907
rect 361488 359864 361540 359873
rect 468024 359864 468076 359916
rect 361672 359703 361724 359712
rect 361672 359669 361681 359703
rect 361681 359669 361715 359703
rect 361715 359669 361724 359703
rect 361672 359660 361724 359669
rect 434904 359660 434956 359712
rect 88340 359363 88392 359372
rect 88340 359329 88349 359363
rect 88349 359329 88383 359363
rect 88383 359329 88392 359363
rect 88340 359320 88392 359329
rect 93492 359252 93544 359304
rect 312544 359116 312596 359168
rect 90640 356779 90692 356788
rect 90640 356745 90649 356779
rect 90649 356745 90683 356779
rect 90683 356745 90692 356779
rect 90640 356736 90692 356745
rect 89260 356668 89312 356720
rect 56692 356600 56744 356652
rect 106372 356600 106424 356652
rect 89260 356575 89312 356584
rect 89260 356541 89269 356575
rect 89269 356541 89303 356575
rect 89303 356541 89312 356575
rect 89260 356532 89312 356541
rect 3792 356056 3844 356108
rect 67088 355988 67140 356040
rect 361580 356031 361632 356040
rect 361580 355997 361589 356031
rect 361589 355997 361623 356031
rect 361623 355997 361632 356031
rect 361580 355988 361632 355997
rect 402428 355988 402480 356040
rect 67548 355852 67600 355904
rect 220544 355852 220596 355904
rect 67548 355308 67600 355360
rect 207020 355308 207072 355360
rect 326988 355308 327040 355360
rect 195244 354356 195296 354408
rect 195428 354356 195480 354408
rect 193680 354220 193732 354272
rect 296076 353812 296128 353864
rect 54024 353744 54076 353796
rect 193588 353379 193640 353388
rect 193588 353345 193597 353379
rect 193597 353345 193631 353379
rect 193631 353345 193640 353379
rect 193588 353336 193640 353345
rect 193680 353379 193732 353388
rect 193680 353345 193689 353379
rect 193689 353345 193723 353379
rect 193723 353345 193732 353379
rect 193680 353336 193732 353345
rect 194600 353447 194652 353456
rect 194600 353413 194609 353447
rect 194609 353413 194643 353447
rect 194643 353413 194652 353447
rect 194600 353404 194652 353413
rect 195428 353379 195480 353388
rect 195428 353345 195437 353379
rect 195437 353345 195471 353379
rect 195471 353345 195480 353379
rect 195428 353336 195480 353345
rect 323584 353336 323636 353388
rect 106188 353268 106240 353320
rect 193864 353311 193916 353320
rect 193864 353277 193873 353311
rect 193873 353277 193907 353311
rect 193907 353277 193916 353311
rect 193864 353268 193916 353277
rect 366364 351636 366416 351688
rect 451464 349503 451516 349512
rect 451464 349469 451473 349503
rect 451473 349469 451507 349503
rect 451507 349469 451516 349503
rect 451464 349460 451516 349469
rect 9404 349324 9456 349376
rect 99840 349052 99892 349104
rect 100668 349052 100720 349104
rect 99840 348508 99892 348560
rect 99656 348440 99708 348492
rect 4620 348279 4672 348288
rect 4620 348245 4629 348279
rect 4629 348245 4663 348279
rect 4663 348245 4672 348279
rect 4620 348236 4672 348245
rect 470600 348372 470652 348424
rect 232320 348304 232372 348356
rect 100944 348236 100996 348288
rect 485412 346851 485464 346860
rect 485412 346817 485421 346851
rect 485421 346817 485455 346851
rect 485455 346817 485464 346851
rect 485412 346808 485464 346817
rect 485596 346851 485648 346860
rect 485596 346817 485605 346851
rect 485605 346817 485639 346851
rect 485639 346817 485648 346851
rect 485596 346808 485648 346817
rect 420920 346604 420972 346656
rect 5264 344428 5316 344480
rect 233332 344267 233384 344276
rect 233332 344233 233341 344267
rect 233341 344233 233375 344267
rect 233375 344233 233384 344267
rect 233332 344224 233384 344233
rect 232688 344131 232740 344140
rect 232688 344097 232697 344131
rect 232697 344097 232731 344131
rect 232731 344097 232740 344131
rect 232688 344088 232740 344097
rect 257068 344088 257120 344140
rect 432604 344020 432656 344072
rect 7932 343884 7984 343936
rect 232964 343927 233016 343936
rect 232964 343893 232973 343927
rect 232973 343893 233007 343927
rect 233007 343893 233016 343927
rect 232964 343884 233016 343893
rect 393228 339668 393280 339720
rect 344744 339235 344796 339244
rect 344744 339201 344753 339235
rect 344753 339201 344787 339235
rect 344787 339201 344796 339235
rect 344744 339192 344796 339201
rect 360384 339192 360436 339244
rect 79784 339124 79836 339176
rect 344928 339031 344980 339040
rect 344928 338997 344937 339031
rect 344937 338997 344971 339031
rect 344971 338997 344980 339031
rect 344928 338988 344980 338997
rect 385132 338147 385184 338156
rect 385132 338113 385141 338147
rect 385141 338113 385175 338147
rect 385175 338113 385184 338147
rect 385132 338104 385184 338113
rect 385224 338147 385276 338156
rect 385224 338113 385233 338147
rect 385233 338113 385267 338147
rect 385267 338113 385276 338147
rect 385224 338104 385276 338113
rect 312268 337696 312320 337748
rect 2964 337492 3016 337544
rect 218704 337535 218756 337544
rect 218704 337501 218713 337535
rect 218713 337501 218747 337535
rect 218747 337501 218756 337535
rect 218704 337492 218756 337501
rect 312360 337492 312412 337544
rect 318800 337492 318852 337544
rect 231032 337424 231084 337476
rect 426900 337424 426952 337476
rect 218520 337399 218572 337408
rect 218520 337365 218529 337399
rect 218529 337365 218563 337399
rect 218563 337365 218572 337399
rect 218520 337356 218572 337365
rect 268752 337356 268804 337408
rect 3148 336676 3200 336728
rect 5356 336676 5408 336728
rect 106188 336064 106240 336116
rect 106372 335971 106424 335980
rect 106372 335937 106381 335971
rect 106381 335937 106415 335971
rect 106415 335937 106424 335971
rect 106372 335928 106424 335937
rect 137928 335860 137980 335912
rect 4068 335724 4120 335776
rect 193588 335724 193640 335776
rect 115940 335316 115992 335368
rect 365812 334679 365864 334688
rect 365812 334645 365821 334679
rect 365821 334645 365855 334679
rect 365855 334645 365864 334679
rect 365812 334636 365864 334645
rect 310612 334364 310664 334416
rect 385224 334296 385276 334348
rect 310612 334271 310664 334280
rect 310612 334237 310621 334271
rect 310621 334237 310655 334271
rect 310655 334237 310664 334271
rect 310612 334228 310664 334237
rect 310796 334271 310848 334280
rect 310796 334237 310805 334271
rect 310805 334237 310839 334271
rect 310839 334237 310848 334271
rect 310796 334228 310848 334237
rect 390928 334228 390980 334280
rect 311072 334160 311124 334212
rect 89076 334092 89128 334144
rect 318156 334024 318208 334076
rect 331772 334160 331824 334212
rect 38844 333208 38896 333260
rect 175556 333140 175608 333192
rect 176016 333072 176068 333124
rect 9128 333004 9180 333056
rect 401140 333004 401192 333056
rect 9128 332800 9180 332852
rect 175740 332800 175792 332852
rect 463700 332596 463752 332648
rect 3608 332528 3660 332580
rect 441988 332528 442040 332580
rect 311256 331372 311308 331424
rect 363512 331211 363564 331220
rect 363512 331177 363521 331211
rect 363521 331177 363555 331211
rect 363555 331177 363564 331211
rect 363512 331168 363564 331177
rect 417516 329740 417568 329792
rect 417792 329740 417844 329792
rect 417884 329536 417936 329588
rect 381452 329443 381504 329452
rect 381452 329409 381461 329443
rect 381461 329409 381495 329443
rect 381495 329409 381504 329443
rect 381452 329400 381504 329409
rect 438308 329443 438360 329452
rect 438308 329409 438317 329443
rect 438317 329409 438351 329443
rect 438351 329409 438360 329443
rect 438308 329400 438360 329409
rect 438492 329443 438544 329452
rect 438492 329409 438501 329443
rect 438501 329409 438535 329443
rect 438535 329409 438544 329443
rect 438492 329400 438544 329409
rect 439964 329332 440016 329384
rect 48228 329264 48280 329316
rect 417516 329264 417568 329316
rect 477684 329264 477736 329316
rect 46204 329196 46256 329248
rect 5264 328992 5316 329044
rect 381452 328992 381504 329044
rect 481732 328992 481784 329044
rect 5172 327700 5224 327752
rect 423772 327360 423824 327412
rect 423956 327267 424008 327276
rect 423956 327233 423965 327267
rect 423965 327233 423999 327267
rect 423999 327233 424008 327267
rect 423956 327224 424008 327233
rect 14464 326612 14516 326664
rect 93308 326179 93360 326188
rect 93308 326145 93317 326179
rect 93317 326145 93351 326179
rect 93351 326145 93360 326179
rect 93308 326136 93360 326145
rect 93492 326179 93544 326188
rect 93492 326145 93501 326179
rect 93501 326145 93535 326179
rect 93535 326145 93544 326179
rect 93492 326136 93544 326145
rect 117780 326136 117832 326188
rect 483020 325932 483072 325984
rect 360844 325728 360896 325780
rect 4712 325524 4764 325576
rect 331588 325091 331640 325100
rect 331588 325057 331597 325091
rect 331597 325057 331631 325091
rect 331631 325057 331640 325091
rect 331588 325048 331640 325057
rect 331772 325091 331824 325100
rect 331772 325057 331781 325091
rect 331781 325057 331815 325091
rect 331815 325057 331824 325091
rect 331772 325048 331824 325057
rect 385224 325048 385276 325100
rect 282276 325023 282328 325032
rect 282276 324989 282285 325023
rect 282285 324989 282319 325023
rect 282319 324989 282328 325023
rect 282276 324980 282328 324989
rect 385040 324980 385092 325032
rect 9220 324844 9272 324896
rect 423864 324844 423916 324896
rect 400036 322872 400088 322924
rect 495440 322872 495492 322924
rect 348424 322711 348476 322720
rect 348424 322677 348433 322711
rect 348433 322677 348467 322711
rect 348467 322677 348476 322711
rect 348424 322668 348476 322677
rect 3608 321580 3660 321632
rect 314476 321580 314528 321632
rect 401508 320152 401560 320204
rect 313832 319404 313884 319456
rect 342260 319107 342312 319116
rect 342260 319073 342269 319107
rect 342269 319073 342303 319107
rect 342303 319073 342312 319107
rect 342260 319064 342312 319073
rect 342536 319064 342588 319116
rect 340972 318860 341024 318912
rect 342076 318860 342128 318912
rect 182088 317407 182140 317416
rect 182088 317373 182097 317407
rect 182097 317373 182131 317407
rect 182131 317373 182140 317407
rect 182088 317364 182140 317373
rect 11704 317228 11756 317280
rect 481824 314347 481876 314356
rect 481824 314313 481833 314347
rect 481833 314313 481867 314347
rect 481867 314313 481876 314347
rect 481824 314304 481876 314313
rect 481732 314211 481784 314220
rect 481732 314177 481741 314211
rect 481741 314177 481775 314211
rect 481775 314177 481784 314211
rect 481732 314168 481784 314177
rect 64788 313216 64840 313268
rect 495440 313216 495492 313268
rect 7564 311856 7616 311908
rect 184480 312103 184532 312112
rect 184480 312069 184498 312103
rect 184498 312069 184532 312103
rect 184480 312060 184532 312069
rect 412364 312060 412416 312112
rect 243084 311924 243136 311976
rect 23388 310700 23440 310752
rect 426716 308728 426768 308780
rect 426992 308728 427044 308780
rect 380900 308592 380952 308644
rect 445760 308660 445812 308712
rect 264612 308524 264664 308576
rect 445760 308388 445812 308440
rect 462320 308388 462372 308440
rect 483020 307776 483072 307828
rect 495440 307776 495492 307828
rect 140780 307096 140832 307148
rect 180800 307096 180852 307148
rect 140780 307003 140832 307012
rect 140780 306969 140789 307003
rect 140789 306969 140823 307003
rect 140823 306969 140832 307003
rect 140780 306960 140832 306969
rect 140872 306935 140924 306944
rect 140872 306901 140881 306935
rect 140881 306901 140915 306935
rect 140915 306901 140924 306935
rect 141240 306935 141292 306944
rect 140872 306892 140924 306901
rect 141240 306901 141249 306935
rect 141249 306901 141283 306935
rect 141283 306901 141292 306935
rect 141240 306892 141292 306901
rect 351184 306348 351236 306400
rect 22100 306187 22152 306196
rect 22100 306153 22109 306187
rect 22109 306153 22143 306187
rect 22143 306153 22152 306187
rect 22100 306144 22152 306153
rect 21640 306051 21692 306060
rect 21640 306017 21649 306051
rect 21649 306017 21683 306051
rect 21683 306017 21692 306051
rect 21640 306008 21692 306017
rect 71872 306008 71924 306060
rect 21548 305804 21600 305856
rect 61108 304852 61160 304904
rect 11428 304784 11480 304836
rect 3884 304716 3936 304768
rect 5816 304716 5868 304768
rect 51448 304759 51500 304768
rect 51448 304725 51457 304759
rect 51457 304725 51491 304759
rect 51491 304725 51500 304759
rect 51448 304716 51500 304725
rect 153384 304716 153436 304768
rect 5908 304512 5960 304564
rect 4712 304215 4764 304224
rect 4712 304181 4721 304215
rect 4721 304181 4755 304215
rect 4755 304181 4764 304215
rect 4712 304172 4764 304181
rect 495624 304172 495676 304224
rect 4160 303084 4212 303136
rect 263600 301588 263652 301640
rect 261116 301495 261168 301504
rect 261116 301461 261125 301495
rect 261125 301461 261159 301495
rect 261159 301461 261168 301495
rect 261116 301452 261168 301461
rect 262312 301452 262364 301504
rect 344744 301452 344796 301504
rect 483756 301452 483808 301504
rect 344744 301112 344796 301164
rect 201960 301044 202012 301096
rect 193864 300908 193916 300960
rect 7840 300092 7892 300144
rect 495440 300092 495492 300144
rect 3884 298324 3936 298376
rect 131120 295944 131172 295996
rect 132408 295944 132460 295996
rect 204996 296148 205048 296200
rect 414388 296191 414440 296200
rect 414388 296157 414397 296191
rect 414397 296157 414431 296191
rect 414431 296157 414440 296191
rect 414388 296148 414440 296157
rect 262312 296012 262364 296064
rect 259092 295808 259144 295860
rect 131120 295740 131172 295792
rect 8300 295604 8352 295656
rect 112168 295715 112220 295724
rect 112168 295681 112176 295715
rect 112176 295681 112210 295715
rect 112210 295681 112220 295715
rect 112536 295715 112588 295724
rect 112168 295672 112220 295681
rect 112536 295681 112545 295715
rect 112545 295681 112579 295715
rect 112579 295681 112588 295715
rect 112536 295672 112588 295681
rect 114468 295672 114520 295724
rect 496268 295672 496320 295724
rect 311072 295604 311124 295656
rect 259460 295536 259512 295588
rect 392124 295468 392176 295520
rect 244372 295264 244424 295316
rect 495440 295264 495492 295316
rect 324964 293972 325016 294024
rect 274732 293335 274784 293344
rect 274732 293301 274741 293335
rect 274741 293301 274775 293335
rect 274775 293301 274784 293335
rect 274732 293292 274784 293301
rect 367100 292884 367152 292936
rect 70584 292408 70636 292460
rect 137928 292383 137980 292392
rect 137928 292349 137937 292383
rect 137937 292349 137971 292383
rect 137971 292349 137980 292383
rect 137928 292340 137980 292349
rect 240140 292204 240192 292256
rect 340880 291363 340932 291372
rect 340880 291329 340889 291363
rect 340889 291329 340923 291363
rect 340923 291329 340932 291363
rect 340880 291320 340932 291329
rect 341432 291363 341484 291372
rect 341432 291329 341441 291363
rect 341441 291329 341475 291363
rect 341475 291329 341484 291363
rect 341432 291320 341484 291329
rect 393320 291320 393372 291372
rect 195060 291184 195112 291236
rect 341340 291252 341392 291304
rect 341248 291184 341300 291236
rect 3608 289824 3660 289876
rect 312452 289824 312504 289876
rect 92940 288099 92992 288108
rect 92940 288065 92949 288099
rect 92949 288065 92983 288099
rect 92983 288065 92992 288099
rect 92940 288056 92992 288065
rect 93124 288099 93176 288108
rect 93124 288065 93133 288099
rect 93133 288065 93167 288099
rect 93167 288065 93176 288099
rect 93124 288056 93176 288065
rect 255688 288056 255740 288108
rect 59636 287852 59688 287904
rect 273628 287011 273680 287020
rect 273628 286977 273637 287011
rect 273637 286977 273671 287011
rect 273671 286977 273680 287011
rect 273628 286968 273680 286977
rect 273812 287011 273864 287020
rect 273812 286977 273821 287011
rect 273821 286977 273855 287011
rect 273855 286977 273864 287011
rect 273812 286968 273864 286977
rect 108304 286900 108356 286952
rect 495440 286900 495492 286952
rect 273996 286875 274048 286884
rect 273996 286841 274005 286875
rect 274005 286841 274039 286875
rect 274039 286841 274048 286875
rect 273996 286832 274048 286841
rect 244464 283883 244516 283892
rect 244464 283849 244473 283883
rect 244473 283849 244507 283883
rect 244507 283849 244516 283883
rect 244464 283840 244516 283849
rect 134340 283704 134392 283756
rect 243084 283679 243136 283688
rect 243084 283645 243093 283679
rect 243093 283645 243127 283679
rect 243127 283645 243136 283679
rect 243084 283636 243136 283645
rect 263600 283704 263652 283756
rect 297640 283704 297692 283756
rect 296904 283636 296956 283688
rect 244464 283500 244516 283552
rect 257160 283500 257212 283552
rect 296076 283339 296128 283348
rect 296076 283305 296085 283339
rect 296085 283305 296119 283339
rect 296119 283305 296128 283339
rect 296076 283296 296128 283305
rect 483020 283339 483072 283348
rect 483020 283305 483029 283339
rect 483029 283305 483063 283339
rect 483063 283305 483072 283339
rect 483020 283296 483072 283305
rect 297640 283203 297692 283212
rect 297640 283169 297649 283203
rect 297649 283169 297683 283203
rect 297683 283169 297692 283203
rect 297640 283160 297692 283169
rect 296720 283135 296772 283144
rect 296720 283101 296729 283135
rect 296729 283101 296763 283135
rect 296763 283101 296772 283135
rect 296720 283092 296772 283101
rect 296904 283024 296956 283076
rect 296720 282752 296772 282804
rect 296076 282659 296128 282668
rect 296076 282625 296085 282659
rect 296085 282625 296119 282659
rect 296119 282625 296128 282659
rect 296076 282616 296128 282625
rect 296904 282659 296956 282668
rect 296904 282625 296913 282659
rect 296913 282625 296947 282659
rect 296947 282625 296956 282659
rect 296904 282616 296956 282625
rect 321468 282548 321520 282600
rect 296076 282480 296128 282532
rect 337752 282140 337804 282192
rect 367560 282140 367612 282192
rect 369216 282004 369268 282056
rect 227904 281528 227956 281580
rect 495440 281528 495492 281580
rect 5632 281324 5684 281376
rect 329748 280483 329800 280492
rect 329748 280449 329757 280483
rect 329757 280449 329791 280483
rect 329791 280449 329800 280483
rect 329748 280440 329800 280449
rect 406292 280440 406344 280492
rect 135904 280236 135956 280288
rect 264612 279463 264664 279472
rect 264612 279429 264646 279463
rect 264646 279429 264664 279463
rect 264612 279420 264664 279429
rect 263600 279352 263652 279404
rect 266360 279352 266412 279404
rect 426900 279148 426952 279200
rect 176936 277899 176988 277908
rect 176936 277865 176945 277899
rect 176945 277865 176979 277899
rect 176979 277865 176988 277899
rect 176936 277856 176988 277865
rect 248696 276131 248748 276140
rect 248696 276097 248705 276131
rect 248705 276097 248739 276131
rect 248739 276097 248748 276131
rect 248696 276088 248748 276097
rect 248604 276063 248656 276072
rect 248604 276029 248613 276063
rect 248613 276029 248647 276063
rect 248647 276029 248656 276063
rect 248604 276020 248656 276029
rect 125876 273912 125928 273964
rect 158904 273955 158956 273964
rect 158904 273921 158912 273955
rect 158912 273921 158946 273955
rect 158946 273921 158956 273955
rect 158904 273912 158956 273921
rect 159088 273955 159140 273964
rect 159088 273921 159097 273955
rect 159097 273921 159131 273955
rect 159131 273921 159140 273955
rect 159088 273912 159140 273921
rect 159272 273955 159324 273964
rect 159272 273921 159281 273955
rect 159281 273921 159315 273955
rect 159315 273921 159324 273955
rect 159272 273912 159324 273921
rect 248236 273912 248288 273964
rect 402796 273912 402848 273964
rect 158996 273887 159048 273896
rect 158996 273853 159005 273887
rect 159005 273853 159039 273887
rect 159039 273853 159048 273887
rect 158996 273844 159048 273853
rect 248604 273844 248656 273896
rect 89168 273708 89220 273760
rect 3240 273300 3292 273352
rect 3608 273164 3660 273216
rect 207112 273164 207164 273216
rect 420552 272663 420604 272672
rect 420552 272629 420561 272663
rect 420561 272629 420595 272663
rect 420595 272629 420604 272663
rect 420552 272620 420604 272629
rect 373080 271328 373132 271380
rect 375472 271328 375524 271380
rect 221464 271124 221516 271176
rect 310704 271124 310756 271176
rect 373080 271167 373132 271176
rect 373080 271133 373089 271167
rect 373089 271133 373123 271167
rect 373123 271133 373132 271167
rect 373080 271124 373132 271133
rect 406384 271056 406436 271108
rect 373816 270827 373868 270836
rect 373816 270793 373825 270827
rect 373825 270793 373859 270827
rect 373859 270793 373868 270827
rect 373816 270784 373868 270793
rect 92296 270283 92348 270292
rect 92296 270249 92305 270283
rect 92305 270249 92339 270283
rect 92339 270249 92348 270283
rect 92296 270240 92348 270249
rect 296076 270036 296128 270088
rect 92296 269900 92348 269952
rect 298836 269900 298888 269952
rect 141240 267860 141292 267912
rect 228916 267903 228968 267912
rect 228916 267869 228925 267903
rect 228925 267869 228959 267903
rect 228959 267869 228968 267903
rect 228916 267860 228968 267869
rect 310244 267860 310296 267912
rect 3608 267724 3660 267776
rect 229100 267767 229152 267776
rect 229100 267733 229109 267767
rect 229109 267733 229143 267767
rect 229143 267733 229152 267767
rect 229100 267724 229152 267733
rect 252560 267724 252612 267776
rect 315488 267724 315540 267776
rect 495440 267724 495492 267776
rect 367284 266815 367336 266824
rect 367284 266781 367293 266815
rect 367293 266781 367327 266815
rect 367327 266781 367336 266815
rect 367284 266772 367336 266781
rect 367468 266815 367520 266824
rect 367468 266781 367477 266815
rect 367477 266781 367511 266815
rect 367511 266781 367520 266815
rect 367468 266772 367520 266781
rect 486976 266815 487028 266824
rect 486976 266781 486985 266815
rect 486985 266781 487019 266815
rect 487019 266781 487028 266815
rect 486976 266772 487028 266781
rect 299388 266704 299440 266756
rect 53932 266636 53984 266688
rect 485596 266679 485648 266688
rect 485596 266645 485605 266679
rect 485605 266645 485639 266679
rect 485639 266645 485648 266679
rect 485596 266636 485648 266645
rect 36360 266339 36412 266348
rect 36360 266305 36369 266339
rect 36369 266305 36403 266339
rect 36403 266305 36412 266339
rect 36360 266296 36412 266305
rect 86868 265752 86920 265804
rect 6736 265684 6788 265736
rect 78128 264163 78180 264172
rect 78128 264129 78162 264163
rect 78162 264129 78180 264163
rect 78128 264120 78180 264129
rect 77852 264095 77904 264104
rect 77852 264061 77861 264095
rect 77861 264061 77895 264095
rect 77895 264061 77904 264095
rect 77852 264052 77904 264061
rect 9036 263916 9088 263968
rect 79232 263959 79284 263968
rect 79232 263925 79241 263959
rect 79241 263925 79275 263959
rect 79275 263925 79284 263959
rect 98736 263959 98788 263968
rect 79232 263916 79284 263925
rect 98736 263925 98745 263959
rect 98745 263925 98779 263959
rect 98779 263925 98788 263959
rect 98736 263916 98788 263925
rect 331404 263916 331456 263968
rect 207204 262556 207256 262608
rect 207020 262420 207072 262472
rect 207388 262463 207440 262472
rect 207388 262429 207397 262463
rect 207397 262429 207431 262463
rect 207431 262429 207440 262463
rect 207388 262420 207440 262429
rect 402980 262420 403032 262472
rect 130476 261264 130528 261316
rect 158812 261264 158864 261316
rect 125784 261196 125836 261248
rect 125876 261035 125928 261044
rect 125876 261001 125893 261035
rect 125893 261001 125927 261035
rect 125927 261001 125928 261035
rect 125876 260992 125928 261001
rect 273812 260992 273864 261044
rect 125324 260899 125376 260908
rect 125324 260865 125333 260899
rect 125333 260865 125367 260899
rect 125367 260865 125376 260899
rect 125324 260856 125376 260865
rect 125784 260899 125836 260908
rect 125784 260865 125787 260899
rect 125787 260865 125836 260899
rect 125784 260856 125836 260865
rect 125876 260856 125928 260908
rect 319812 260924 319864 260976
rect 131580 260856 131632 260908
rect 319904 260856 319956 260908
rect 339960 260244 340012 260296
rect 317696 260151 317748 260160
rect 317696 260117 317705 260151
rect 317705 260117 317739 260151
rect 317739 260117 317748 260151
rect 317696 260108 317748 260117
rect 331220 260108 331272 260160
rect 180800 259224 180852 259276
rect 180984 259224 181036 259276
rect 232688 259224 232740 259276
rect 268384 259156 268436 259208
rect 180892 259131 180944 259140
rect 180892 259097 180901 259131
rect 180901 259097 180935 259131
rect 180935 259097 180944 259131
rect 180892 259088 180944 259097
rect 180800 259063 180852 259072
rect 180800 259029 180809 259063
rect 180809 259029 180843 259063
rect 180843 259029 180852 259063
rect 181260 259063 181312 259072
rect 180800 259020 180852 259029
rect 181260 259029 181269 259063
rect 181269 259029 181303 259063
rect 181303 259029 181312 259063
rect 181260 259020 181312 259029
rect 347044 258068 347096 258120
rect 495440 258068 495492 258120
rect 483756 257635 483808 257644
rect 483756 257601 483765 257635
rect 483765 257601 483799 257635
rect 483799 257601 483808 257635
rect 483756 257592 483808 257601
rect 181260 257524 181312 257576
rect 321928 257388 321980 257440
rect 470508 257023 470560 257032
rect 470508 256989 470517 257023
rect 470517 256989 470551 257023
rect 470551 256989 470560 257023
rect 470508 256980 470560 256989
rect 470600 256887 470652 256896
rect 470600 256853 470609 256887
rect 470609 256853 470643 256887
rect 470643 256853 470652 256887
rect 470600 256844 470652 256853
rect 299388 256683 299440 256692
rect 299388 256649 299397 256683
rect 299397 256649 299431 256683
rect 299431 256649 299440 256683
rect 299388 256640 299440 256649
rect 299204 256547 299256 256556
rect 299204 256513 299213 256547
rect 299213 256513 299247 256547
rect 299247 256513 299256 256547
rect 299204 256504 299256 256513
rect 485596 256504 485648 256556
rect 298836 256479 298888 256488
rect 298836 256445 298845 256479
rect 298845 256445 298879 256479
rect 298879 256445 298888 256479
rect 298836 256436 298888 256445
rect 333980 256436 334032 256488
rect 334348 256436 334400 256488
rect 310428 256368 310480 256420
rect 117596 256300 117648 256352
rect 333980 256028 334032 256080
rect 371148 256028 371200 256080
rect 310060 255960 310112 256012
rect 310428 255960 310480 256012
rect 334072 255960 334124 256012
rect 371424 255960 371476 256012
rect 263784 255212 263836 255264
rect 381452 255212 381504 255264
rect 220544 254915 220596 254924
rect 220544 254881 220553 254915
rect 220553 254881 220587 254915
rect 220587 254881 220596 254915
rect 220544 254872 220596 254881
rect 396632 254847 396684 254856
rect 396632 254813 396641 254847
rect 396641 254813 396675 254847
rect 396675 254813 396684 254847
rect 396632 254804 396684 254813
rect 219808 254736 219860 254788
rect 219256 254668 219308 254720
rect 263784 254668 263836 254720
rect 349068 254124 349120 254176
rect 117596 252875 117648 252884
rect 117596 252841 117605 252875
rect 117605 252841 117639 252875
rect 117639 252841 117648 252875
rect 117596 252832 117648 252841
rect 3240 252696 3292 252748
rect 9312 252628 9364 252680
rect 117780 252671 117832 252680
rect 117780 252637 117789 252671
rect 117789 252637 117823 252671
rect 117823 252637 117832 252671
rect 117780 252628 117832 252637
rect 414664 252628 414716 252680
rect 260656 252560 260708 252612
rect 444012 252195 444064 252204
rect 444012 252161 444021 252195
rect 444021 252161 444055 252195
rect 444055 252161 444064 252195
rect 444012 252152 444064 252161
rect 444104 252127 444156 252136
rect 444104 252093 444113 252127
rect 444113 252093 444147 252127
rect 444147 252093 444156 252127
rect 444104 252084 444156 252093
rect 444196 252127 444248 252136
rect 444196 252093 444205 252127
rect 444205 252093 444239 252127
rect 444239 252093 444248 252127
rect 444196 252084 444248 252093
rect 336096 251948 336148 252000
rect 274732 251132 274784 251184
rect 495440 251132 495492 251184
rect 4620 251064 4672 251116
rect 266360 251064 266412 251116
rect 232320 250971 232372 250980
rect 232320 250937 232329 250971
rect 232329 250937 232363 250971
rect 232363 250937 232372 250971
rect 232320 250928 232372 250937
rect 254216 250860 254268 250912
rect 257252 250860 257304 250912
rect 303160 250019 303212 250028
rect 303160 249985 303169 250019
rect 303169 249985 303203 250019
rect 303203 249985 303212 250019
rect 303160 249976 303212 249985
rect 361580 249976 361632 250028
rect 12992 249772 13044 249824
rect 315120 248727 315172 248736
rect 315120 248693 315129 248727
rect 315129 248693 315163 248727
rect 315163 248693 315172 248727
rect 315120 248684 315172 248693
rect 311440 244332 311492 244384
rect 315764 240907 315816 240916
rect 315764 240873 315773 240907
rect 315773 240873 315807 240907
rect 315807 240873 315816 240907
rect 315764 240864 315816 240873
rect 468024 240907 468076 240916
rect 468024 240873 468033 240907
rect 468033 240873 468067 240907
rect 468067 240873 468076 240907
rect 468024 240864 468076 240873
rect 467380 240635 467432 240644
rect 467380 240601 467389 240635
rect 467389 240601 467423 240635
rect 467423 240601 467432 240635
rect 467380 240592 467432 240601
rect 467840 240635 467892 240644
rect 467840 240601 467849 240635
rect 467849 240601 467883 240635
rect 467883 240601 467892 240635
rect 467840 240592 467892 240601
rect 496268 240592 496320 240644
rect 467656 240567 467708 240576
rect 467656 240533 467665 240567
rect 467665 240533 467699 240567
rect 467699 240533 467708 240567
rect 467656 240524 467708 240533
rect 467748 240567 467800 240576
rect 467748 240533 467757 240567
rect 467757 240533 467791 240567
rect 467791 240533 467800 240567
rect 467748 240524 467800 240533
rect 372620 238484 372672 238536
rect 373080 238484 373132 238536
rect 20536 237575 20588 237584
rect 20536 237541 20545 237575
rect 20545 237541 20579 237575
rect 20579 237541 20588 237575
rect 430948 237575 431000 237584
rect 20536 237532 20588 237541
rect 430948 237541 430957 237575
rect 430957 237541 430991 237575
rect 430991 237541 431000 237575
rect 430948 237532 431000 237541
rect 59452 237464 59504 237516
rect 372620 237396 372672 237448
rect 430764 237439 430816 237448
rect 430764 237405 430773 237439
rect 430773 237405 430807 237439
rect 430807 237405 430816 237439
rect 430764 237396 430816 237405
rect 430948 237396 431000 237448
rect 435272 237396 435324 237448
rect 77852 236648 77904 236700
rect 133236 236648 133288 236700
rect 5172 236308 5224 236360
rect 61108 236351 61160 236360
rect 61108 236317 61117 236351
rect 61117 236317 61151 236351
rect 61151 236317 61160 236351
rect 61108 236308 61160 236317
rect 77852 236308 77904 236360
rect 342536 236351 342588 236360
rect 342536 236317 342545 236351
rect 342545 236317 342579 236351
rect 342579 236317 342588 236351
rect 342536 236308 342588 236317
rect 416136 236308 416188 236360
rect 61476 236240 61528 236292
rect 62488 236215 62540 236224
rect 62488 236181 62497 236215
rect 62497 236181 62531 236215
rect 62531 236181 62540 236215
rect 62488 236172 62540 236181
rect 155960 236172 156012 236224
rect 341156 236215 341208 236224
rect 341156 236181 341165 236215
rect 341165 236181 341199 236215
rect 341199 236181 341208 236215
rect 341156 236172 341208 236181
rect 342352 236172 342404 236224
rect 240324 232475 240376 232484
rect 240324 232441 240333 232475
rect 240333 232441 240367 232475
rect 240367 232441 240376 232475
rect 240324 232432 240376 232441
rect 216220 231523 216272 231532
rect 216220 231489 216229 231523
rect 216229 231489 216263 231523
rect 216263 231489 216272 231523
rect 216220 231480 216272 231489
rect 204352 230800 204404 230852
rect 419080 230979 419132 230988
rect 419080 230945 419089 230979
rect 419089 230945 419123 230979
rect 419123 230945 419132 230979
rect 419080 230936 419132 230945
rect 444196 230936 444248 230988
rect 126980 230732 127032 230784
rect 418712 230732 418764 230784
rect 153384 229823 153436 229832
rect 153384 229789 153393 229823
rect 153393 229789 153427 229823
rect 153427 229789 153436 229823
rect 153384 229780 153436 229789
rect 153476 229823 153528 229832
rect 153476 229789 153485 229823
rect 153485 229789 153519 229823
rect 153519 229789 153528 229823
rect 153476 229780 153528 229789
rect 167828 228395 167880 228404
rect 167828 228361 167837 228395
rect 167837 228361 167871 228395
rect 167871 228361 167880 228395
rect 167828 228352 167880 228361
rect 167460 228259 167512 228268
rect 167460 228225 167469 228259
rect 167469 228225 167503 228259
rect 167503 228225 167512 228259
rect 167460 228216 167512 228225
rect 167184 228191 167236 228200
rect 167184 228157 167193 228191
rect 167193 228157 167227 228191
rect 167227 228157 167236 228191
rect 167184 228148 167236 228157
rect 167368 228191 167420 228200
rect 167368 228157 167377 228191
rect 167377 228157 167411 228191
rect 167411 228157 167420 228191
rect 167368 228148 167420 228157
rect 175832 228148 175884 228200
rect 180800 228148 180852 228200
rect 315580 228012 315632 228064
rect 137192 227715 137244 227724
rect 137192 227681 137201 227715
rect 137201 227681 137235 227715
rect 137235 227681 137244 227715
rect 137192 227672 137244 227681
rect 167644 227672 167696 227724
rect 329748 227672 329800 227724
rect 137192 227536 137244 227588
rect 135628 227171 135680 227180
rect 135628 227137 135637 227171
rect 135637 227137 135671 227171
rect 135671 227137 135680 227171
rect 135628 227128 135680 227137
rect 135904 227171 135956 227180
rect 135904 227137 135913 227171
rect 135913 227137 135947 227171
rect 135947 227137 135956 227171
rect 135904 227128 135956 227137
rect 135996 227171 136048 227180
rect 135996 227137 136006 227171
rect 136006 227137 136040 227171
rect 136040 227137 136048 227171
rect 135996 227128 136048 227137
rect 136548 227060 136600 227112
rect 175648 227196 175700 227248
rect 137192 227103 137244 227112
rect 137192 227069 137201 227103
rect 137201 227069 137235 227103
rect 137235 227069 137244 227103
rect 137192 227060 137244 227069
rect 167644 227060 167696 227112
rect 40592 226924 40644 226976
rect 347044 225675 347096 225684
rect 347044 225641 347053 225675
rect 347053 225641 347087 225675
rect 347087 225641 347096 225675
rect 347044 225632 347096 225641
rect 290280 224995 290332 225004
rect 290280 224961 290289 224995
rect 290289 224961 290323 224995
rect 290323 224961 290332 224995
rect 290280 224952 290332 224961
rect 335912 224952 335964 225004
rect 289820 224791 289872 224800
rect 289820 224757 289829 224791
rect 289829 224757 289863 224791
rect 289863 224757 289872 224791
rect 289820 224748 289872 224757
rect 100852 224587 100904 224596
rect 100852 224553 100861 224587
rect 100861 224553 100895 224587
rect 100895 224553 100904 224587
rect 100852 224544 100904 224553
rect 290004 224587 290056 224596
rect 290004 224553 290013 224587
rect 290013 224553 290047 224587
rect 290047 224553 290056 224587
rect 290004 224544 290056 224553
rect 289820 224408 289872 224460
rect 100944 224383 100996 224392
rect 100944 224349 100953 224383
rect 100953 224349 100987 224383
rect 100987 224349 100996 224383
rect 100944 224340 100996 224349
rect 310796 224340 310848 224392
rect 32772 224204 32824 224256
rect 289636 224247 289688 224256
rect 289636 224213 289645 224247
rect 289645 224213 289679 224247
rect 289679 224213 289688 224247
rect 289636 224204 289688 224213
rect 3056 223728 3108 223780
rect 5908 223728 5960 223780
rect 126980 223524 127032 223576
rect 127532 223524 127584 223576
rect 141424 223524 141476 223576
rect 142068 223524 142120 223576
rect 134524 223456 134576 223508
rect 228088 223524 228140 223576
rect 260840 223524 260892 223576
rect 467656 223456 467708 223508
rect 207388 223388 207440 223440
rect 379520 223388 379572 223440
rect 42064 223320 42116 223372
rect 239036 223320 239088 223372
rect 187608 223252 187660 223304
rect 260472 223295 260524 223304
rect 260472 223261 260481 223295
rect 260481 223261 260515 223295
rect 260515 223261 260524 223295
rect 260472 223252 260524 223261
rect 260564 223252 260616 223304
rect 367284 223320 367336 223372
rect 430580 223252 430632 223304
rect 194416 223184 194468 223236
rect 255964 223184 256016 223236
rect 260748 223184 260800 223236
rect 496636 223184 496688 223236
rect 61844 223116 61896 223168
rect 260564 223116 260616 223168
rect 260656 223159 260708 223168
rect 260656 223125 260665 223159
rect 260665 223125 260699 223159
rect 260699 223125 260708 223159
rect 260656 223116 260708 223125
rect 382280 223116 382332 223168
rect 93676 223048 93728 223100
rect 147772 223048 147824 223100
rect 112260 222980 112312 223032
rect 200396 222980 200448 223032
rect 280528 222980 280580 223032
rect 328460 222980 328512 223032
rect 35164 222912 35216 222964
rect 426808 222912 426860 222964
rect 95056 222844 95108 222896
rect 496360 222844 496412 222896
rect 81808 222776 81860 222828
rect 82728 222776 82780 222828
rect 140872 222776 140924 222828
rect 247132 222776 247184 222828
rect 199936 222708 199988 222760
rect 299756 222708 299808 222760
rect 53840 222640 53892 222692
rect 54668 222640 54720 222692
rect 153200 222640 153252 222692
rect 154028 222640 154080 222692
rect 205824 222640 205876 222692
rect 286508 222640 286560 222692
rect 101404 222572 101456 222624
rect 438492 222572 438544 222624
rect 252560 222504 252612 222556
rect 253388 222504 253440 222556
rect 68560 222368 68612 222420
rect 259184 222368 259236 222420
rect 260656 222368 260708 222420
rect 475384 222368 475436 222420
rect 227536 222300 227588 222352
rect 496728 222300 496780 222352
rect 7196 222232 7248 222284
rect 21640 222232 21692 222284
rect 48688 222232 48740 222284
rect 381084 222232 381136 222284
rect 15568 222164 15620 222216
rect 362224 222164 362276 222216
rect 79784 220779 79836 220788
rect 79784 220745 79793 220779
rect 79793 220745 79827 220779
rect 79827 220745 79836 220779
rect 79784 220736 79836 220745
rect 97080 220779 97132 220788
rect 97080 220745 97089 220779
rect 97089 220745 97123 220779
rect 97123 220745 97132 220779
rect 97080 220736 97132 220745
rect 123392 220779 123444 220788
rect 123392 220745 123401 220779
rect 123401 220745 123435 220779
rect 123435 220745 123444 220779
rect 123392 220736 123444 220745
rect 112536 220668 112588 220720
rect 159088 220668 159140 220720
rect 204996 220736 205048 220788
rect 205456 220736 205508 220788
rect 205640 220779 205692 220788
rect 205640 220745 205649 220779
rect 205649 220745 205683 220779
rect 205683 220745 205692 220779
rect 205640 220736 205692 220745
rect 205732 220736 205784 220788
rect 209044 220736 209096 220788
rect 341248 220736 341300 220788
rect 248696 220668 248748 220720
rect 249708 220668 249760 220720
rect 79416 220643 79468 220652
rect 79416 220609 79425 220643
rect 79425 220609 79459 220643
rect 79459 220609 79468 220643
rect 79416 220600 79468 220609
rect 107660 220600 107712 220652
rect 178316 220643 178368 220652
rect 178316 220609 178325 220643
rect 178325 220609 178359 220643
rect 178359 220609 178368 220643
rect 178316 220600 178368 220609
rect 204996 220643 205048 220652
rect 204996 220609 205005 220643
rect 205005 220609 205039 220643
rect 205039 220609 205048 220643
rect 204996 220600 205048 220609
rect 205180 220643 205232 220652
rect 205180 220609 205188 220643
rect 205188 220609 205222 220643
rect 205222 220609 205232 220643
rect 205180 220600 205232 220609
rect 205272 220643 205324 220652
rect 205272 220609 205281 220643
rect 205281 220609 205315 220643
rect 205315 220609 205324 220643
rect 205272 220600 205324 220609
rect 79324 220575 79376 220584
rect 79324 220541 79333 220575
rect 79333 220541 79367 220575
rect 79367 220541 79376 220575
rect 79324 220532 79376 220541
rect 96620 220575 96672 220584
rect 96620 220541 96629 220575
rect 96629 220541 96663 220575
rect 96663 220541 96672 220575
rect 96620 220532 96672 220541
rect 133236 220575 133288 220584
rect 133236 220541 133245 220575
rect 133245 220541 133279 220575
rect 133279 220541 133288 220575
rect 162768 220575 162820 220584
rect 133236 220532 133288 220541
rect 55036 220507 55088 220516
rect 55036 220473 55045 220507
rect 55045 220473 55079 220507
rect 55079 220473 55088 220507
rect 55036 220464 55088 220473
rect 125784 220464 125836 220516
rect 137928 220464 137980 220516
rect 162768 220541 162777 220575
rect 162777 220541 162811 220575
rect 162811 220541 162820 220575
rect 162768 220532 162820 220541
rect 205364 220575 205416 220584
rect 205364 220541 205373 220575
rect 205373 220541 205407 220575
rect 205407 220541 205416 220575
rect 205364 220532 205416 220541
rect 235264 220643 235316 220652
rect 235264 220609 235273 220643
rect 235273 220609 235307 220643
rect 235307 220609 235316 220643
rect 235264 220600 235316 220609
rect 258908 220668 258960 220720
rect 259276 220711 259328 220720
rect 259276 220677 259285 220711
rect 259285 220677 259319 220711
rect 259319 220677 259328 220711
rect 259276 220668 259328 220677
rect 266084 220668 266136 220720
rect 430948 220668 431000 220720
rect 257436 220643 257488 220652
rect 257436 220609 257445 220643
rect 257445 220609 257479 220643
rect 257479 220609 257488 220643
rect 257436 220600 257488 220609
rect 259092 220643 259144 220652
rect 259092 220609 259096 220643
rect 259096 220609 259130 220643
rect 259130 220609 259144 220643
rect 259092 220600 259144 220609
rect 259184 220643 259236 220652
rect 259184 220609 259193 220643
rect 259193 220609 259227 220643
rect 259227 220609 259236 220643
rect 259460 220643 259512 220652
rect 259184 220600 259236 220609
rect 259460 220609 259468 220643
rect 259468 220609 259502 220643
rect 259502 220609 259512 220643
rect 259460 220600 259512 220609
rect 259644 220600 259696 220652
rect 257160 220575 257212 220584
rect 257160 220541 257169 220575
rect 257169 220541 257203 220575
rect 257203 220541 257212 220575
rect 257160 220532 257212 220541
rect 257252 220575 257304 220584
rect 257252 220541 257261 220575
rect 257261 220541 257295 220575
rect 257295 220541 257304 220575
rect 257252 220532 257304 220541
rect 205548 220464 205600 220516
rect 257344 220464 257396 220516
rect 49976 220439 50028 220448
rect 49976 220405 49985 220439
rect 49985 220405 50019 220439
rect 50019 220405 50028 220439
rect 49976 220396 50028 220405
rect 77760 220439 77812 220448
rect 77760 220405 77769 220439
rect 77769 220405 77803 220439
rect 77803 220405 77812 220439
rect 77760 220396 77812 220405
rect 125324 220192 125376 220244
rect 205272 220396 205324 220448
rect 213184 220396 213236 220448
rect 266636 220532 266688 220584
rect 282920 220600 282972 220652
rect 342536 220532 342588 220584
rect 257620 220464 257672 220516
rect 257712 220439 257764 220448
rect 257712 220405 257721 220439
rect 257721 220405 257755 220439
rect 257755 220405 257764 220439
rect 257712 220396 257764 220405
rect 265072 220439 265124 220448
rect 265072 220405 265081 220439
rect 265081 220405 265115 220439
rect 265115 220405 265124 220439
rect 265072 220396 265124 220405
rect 318524 220464 318576 220516
rect 266544 220396 266596 220448
rect 341340 220396 341392 220448
rect 266636 220328 266688 220380
rect 317236 220192 317288 220244
rect 315672 220124 315724 220176
rect 318708 220124 318760 220176
rect 361672 220124 361724 220176
rect 23020 220056 23072 220108
rect 238484 220056 238536 220108
rect 259644 220056 259696 220108
rect 340420 220056 340472 220108
rect 310612 219988 310664 220040
rect 167184 219920 167236 219972
rect 318340 219920 318392 219972
rect 259460 219852 259512 219904
rect 318708 219852 318760 219904
rect 264980 219784 265032 219836
rect 265072 219784 265124 219836
rect 313188 219784 313240 219836
rect 249708 219716 249760 219768
rect 310336 219716 310388 219768
rect 162768 219648 162820 219700
rect 259092 219648 259144 219700
rect 282920 219648 282972 219700
rect 317144 219648 317196 219700
rect 205180 219580 205232 219632
rect 495992 219580 496044 219632
rect 11796 219555 11848 219564
rect 11796 219521 11805 219555
rect 11805 219521 11839 219555
rect 11839 219521 11848 219555
rect 11796 219512 11848 219521
rect 12808 219555 12860 219564
rect 12808 219521 12817 219555
rect 12817 219521 12851 219555
rect 12851 219521 12860 219555
rect 12808 219512 12860 219521
rect 16212 219555 16264 219564
rect 16212 219521 16221 219555
rect 16221 219521 16255 219555
rect 16255 219521 16264 219555
rect 16212 219512 16264 219521
rect 17224 219555 17276 219564
rect 17224 219521 17233 219555
rect 17233 219521 17267 219555
rect 17267 219521 17276 219555
rect 17224 219512 17276 219521
rect 96068 219555 96120 219564
rect 4436 219444 4488 219496
rect 53748 219487 53800 219496
rect 53748 219453 53757 219487
rect 53757 219453 53791 219487
rect 53791 219453 53800 219487
rect 53748 219444 53800 219453
rect 96068 219521 96077 219555
rect 96077 219521 96111 219555
rect 96111 219521 96120 219555
rect 96068 219512 96120 219521
rect 257160 219512 257212 219564
rect 318432 219512 318484 219564
rect 3608 219376 3660 219428
rect 130384 219376 130436 219428
rect 7840 219308 7892 219360
rect 20536 219308 20588 219360
rect 21548 219308 21600 219360
rect 22928 219351 22980 219360
rect 22928 219317 22937 219351
rect 22937 219317 22971 219351
rect 22971 219317 22980 219351
rect 22928 219308 22980 219317
rect 7748 219240 7800 219292
rect 8484 219172 8536 219224
rect 55496 219308 55548 219360
rect 78128 219351 78180 219360
rect 78128 219317 78137 219351
rect 78137 219317 78171 219351
rect 78171 219317 78180 219351
rect 78128 219308 78180 219317
rect 8208 219104 8260 219156
rect 101496 219308 101548 219360
rect 112996 219308 113048 219360
rect 114376 219351 114428 219360
rect 114376 219317 114385 219351
rect 114385 219317 114419 219351
rect 114419 219317 114428 219351
rect 114376 219308 114428 219317
rect 218520 219308 218572 219360
rect 232964 219351 233016 219360
rect 5448 218968 5500 219020
rect 4620 218900 4672 218952
rect 232964 219317 232973 219351
rect 232973 219317 233007 219351
rect 233007 219317 233016 219351
rect 232964 219308 233016 219317
rect 248328 219351 248380 219360
rect 248328 219317 248337 219351
rect 248337 219317 248371 219351
rect 248371 219317 248380 219351
rect 248328 219308 248380 219317
rect 249432 219308 249484 219360
rect 260748 219308 260800 219360
rect 310980 219036 311032 219088
rect 311532 218968 311584 219020
rect 311808 218900 311860 218952
rect 8576 218832 8628 218884
rect 310796 218832 310848 218884
rect 8760 218764 8812 218816
rect 483848 218764 483900 218816
rect 9496 218696 9548 218748
rect 310888 218696 310940 218748
rect 6920 218628 6972 218680
rect 6736 218560 6788 218612
rect 5724 218492 5776 218544
rect 7288 218424 7340 218476
rect 399484 218016 399536 218068
rect 495440 218016 495492 218068
rect 9496 217719 9548 217728
rect 9496 217685 9505 217719
rect 9505 217685 9539 217719
rect 9539 217685 9548 217719
rect 9496 217676 9548 217685
rect 3608 217608 3660 217660
rect 310520 217608 310572 217660
rect 8392 217540 8444 217592
rect 485412 217540 485464 217592
rect 7472 217472 7524 217524
rect 496360 217472 496412 217524
rect 312544 216792 312596 216844
rect 371148 216928 371200 216980
rect 313188 216724 313240 216776
rect 371148 216767 371200 216776
rect 371148 216733 371157 216767
rect 371157 216733 371191 216767
rect 371191 216733 371200 216767
rect 371148 216724 371200 216733
rect 371424 216767 371476 216776
rect 371424 216733 371433 216767
rect 371433 216733 371467 216767
rect 371467 216733 371476 216767
rect 371424 216724 371476 216733
rect 428924 216860 428976 216912
rect 340420 216656 340472 216708
rect 310520 210400 310572 210452
rect 6000 209516 6052 209568
rect 2872 205980 2924 206032
rect 5632 205980 5684 206032
rect 8668 203872 8720 203924
rect 9496 203915 9548 203924
rect 9496 203881 9505 203915
rect 9505 203881 9539 203915
rect 9539 203881 9548 203915
rect 9496 203872 9548 203881
rect 5632 203668 5684 203720
rect 331220 202784 331272 202836
rect 467380 202784 467432 202836
rect 311072 202104 311124 202156
rect 311808 201968 311860 202020
rect 331220 201900 331272 201952
rect 313832 201424 313884 201476
rect 495440 201424 495492 201476
rect 322204 200812 322256 200864
rect 483848 199971 483900 199980
rect 483848 199937 483857 199971
rect 483857 199937 483891 199971
rect 483891 199937 483900 199971
rect 483848 199928 483900 199937
rect 3240 197752 3292 197804
rect 7564 197752 7616 197804
rect 405924 197276 405976 197328
rect 495440 197276 495492 197328
rect 349804 195372 349856 195424
rect 315764 194964 315816 195016
rect 472624 191836 472676 191888
rect 495440 191836 495492 191888
rect 349804 187688 349856 187740
rect 495440 187688 495492 187740
rect 310336 183948 310388 184000
rect 310336 183651 310388 183660
rect 310336 183617 310344 183651
rect 310344 183617 310378 183651
rect 310378 183617 310388 183651
rect 310336 183608 310388 183617
rect 311624 183744 311676 183796
rect 310796 183676 310848 183728
rect 469864 183676 469916 183728
rect 310704 183651 310756 183660
rect 310704 183617 310713 183651
rect 310713 183617 310747 183651
rect 310747 183617 310756 183651
rect 310704 183608 310756 183617
rect 311808 183608 311860 183660
rect 310612 183540 310664 183592
rect 453028 183540 453080 183592
rect 3056 183404 3108 183456
rect 6092 183404 6144 183456
rect 406384 179775 406436 179784
rect 406384 179741 406393 179775
rect 406393 179741 406427 179775
rect 406427 179741 406436 179775
rect 406384 179732 406436 179741
rect 407396 179639 407448 179648
rect 407396 179605 407405 179639
rect 407405 179605 407439 179639
rect 407439 179605 407448 179639
rect 407396 179596 407448 179605
rect 3332 178848 3384 178900
rect 3976 178848 4028 178900
rect 310704 178508 310756 178560
rect 346860 178508 346912 178560
rect 310888 178304 310940 178356
rect 310520 178236 310572 178288
rect 311532 178236 311584 178288
rect 310428 178211 310480 178220
rect 310428 178177 310437 178211
rect 310437 178177 310471 178211
rect 310471 178177 310480 178211
rect 310428 178168 310480 178177
rect 407396 178168 407448 178220
rect 310704 178143 310756 178152
rect 310704 178109 310713 178143
rect 310713 178109 310747 178143
rect 310747 178109 310756 178143
rect 310704 178100 310756 178109
rect 310796 178032 310848 178084
rect 310244 176171 310296 176180
rect 310244 176137 310253 176171
rect 310253 176137 310287 176171
rect 310287 176137 310296 176171
rect 310244 176128 310296 176137
rect 336188 176171 336240 176180
rect 336188 176137 336197 176171
rect 336197 176137 336231 176171
rect 336231 176137 336240 176171
rect 336188 176128 336240 176137
rect 336556 176171 336608 176180
rect 336556 176137 336565 176171
rect 336565 176137 336599 176171
rect 336599 176137 336608 176171
rect 336556 176128 336608 176137
rect 336096 176103 336148 176112
rect 336096 176069 336105 176103
rect 336105 176069 336139 176103
rect 336139 176069 336148 176103
rect 336096 176060 336148 176069
rect 310704 175992 310756 176044
rect 310980 175992 311032 176044
rect 335912 175967 335964 175976
rect 335912 175933 335921 175967
rect 335921 175933 335955 175967
rect 335955 175933 335964 175967
rect 335912 175924 335964 175933
rect 337476 175831 337528 175840
rect 337476 175797 337485 175831
rect 337485 175797 337519 175831
rect 337519 175797 337528 175831
rect 337476 175788 337528 175797
rect 310244 175584 310296 175636
rect 419540 175584 419592 175636
rect 324964 175176 325016 175228
rect 495440 175176 495492 175228
rect 3332 170144 3384 170196
rect 5172 170008 5224 170060
rect 5080 169940 5132 169992
rect 3976 169804 4028 169856
rect 7380 169804 7432 169856
rect 380624 161984 380676 162036
rect 381084 162027 381136 162036
rect 381084 161993 381093 162027
rect 381093 161993 381127 162027
rect 381127 161993 381136 162027
rect 381084 161984 381136 161993
rect 378784 161916 378836 161968
rect 424048 161984 424100 162036
rect 470508 161916 470560 161968
rect 385040 161891 385092 161900
rect 385040 161857 385049 161891
rect 385049 161857 385083 161891
rect 385083 161857 385092 161891
rect 385040 161848 385092 161857
rect 385224 161891 385276 161900
rect 385224 161857 385233 161891
rect 385233 161857 385267 161891
rect 385267 161857 385276 161891
rect 385224 161848 385276 161857
rect 385592 161891 385644 161900
rect 385592 161857 385601 161891
rect 385601 161857 385635 161891
rect 385635 161857 385644 161891
rect 385592 161848 385644 161857
rect 385776 161891 385828 161900
rect 385776 161857 385785 161891
rect 385785 161857 385819 161891
rect 385819 161857 385828 161891
rect 385776 161848 385828 161857
rect 380164 161780 380216 161832
rect 382188 161780 382240 161832
rect 419080 161848 419132 161900
rect 414848 161687 414900 161696
rect 414848 161653 414857 161687
rect 414857 161653 414891 161687
rect 414891 161653 414900 161687
rect 414848 161644 414900 161653
rect 315948 161440 316000 161492
rect 3332 161100 3384 161152
rect 6460 161100 6512 161152
rect 9128 157088 9180 157140
rect 484216 157131 484268 157140
rect 484216 157097 484225 157131
rect 484225 157097 484259 157131
rect 484259 157097 484268 157131
rect 484216 157088 484268 157097
rect 3148 157020 3200 157072
rect 6368 157020 6420 157072
rect 8944 156884 8996 156936
rect 321468 152643 321520 152652
rect 321468 152609 321477 152643
rect 321477 152609 321511 152643
rect 321511 152609 321520 152643
rect 321468 152600 321520 152609
rect 323584 152643 323636 152652
rect 323584 152609 323593 152643
rect 323593 152609 323627 152643
rect 323627 152609 323636 152643
rect 323584 152600 323636 152609
rect 429200 152532 429252 152584
rect 425704 152056 425756 152108
rect 321928 152031 321980 152040
rect 321928 151997 321937 152031
rect 321937 151997 321971 152031
rect 321971 151997 321980 152031
rect 321928 151988 321980 151997
rect 321652 151920 321704 151972
rect 417516 151988 417568 152040
rect 321376 151852 321428 151904
rect 357348 148223 357400 148232
rect 357348 148189 357357 148223
rect 357357 148189 357391 148223
rect 357391 148189 357400 148223
rect 357348 148180 357400 148189
rect 315212 147500 315264 147552
rect 486976 146888 487028 146940
rect 495532 146888 495584 146940
rect 418160 143488 418212 143540
rect 418804 143488 418856 143540
rect 495440 143488 495492 143540
rect 389364 143191 389416 143200
rect 389364 143157 389373 143191
rect 389373 143157 389407 143191
rect 389407 143157 389416 143191
rect 389364 143148 389416 143157
rect 316592 142808 316644 142860
rect 418160 142808 418212 142860
rect 361488 142740 361540 142792
rect 9772 142307 9824 142316
rect 9772 142273 9781 142307
rect 9781 142273 9815 142307
rect 9815 142273 9824 142307
rect 9772 142264 9824 142273
rect 9772 142128 9824 142180
rect 313832 142128 313884 142180
rect 416136 140607 416188 140616
rect 416136 140573 416145 140607
rect 416145 140573 416179 140607
rect 416179 140573 416188 140607
rect 416136 140564 416188 140573
rect 451648 140564 451700 140616
rect 416412 140539 416464 140548
rect 416412 140505 416446 140539
rect 416446 140505 416464 140539
rect 416412 140496 416464 140505
rect 417424 140428 417476 140480
rect 473636 140428 473688 140480
rect 3332 138932 3384 138984
rect 6552 138932 6604 138984
rect 8392 136416 8444 136468
rect 9128 136416 9180 136468
rect 8484 136212 8536 136264
rect 8944 136212 8996 136264
rect 8576 133084 8628 133136
rect 9036 133016 9088 133068
rect 9220 133059 9272 133068
rect 9220 133025 9229 133059
rect 9229 133025 9263 133059
rect 9263 133025 9272 133059
rect 9220 133016 9272 133025
rect 9404 133016 9456 133068
rect 9496 132991 9548 133000
rect 9496 132957 9505 132991
rect 9505 132957 9539 132991
rect 9539 132957 9548 132991
rect 9496 132948 9548 132957
rect 369308 132948 369360 133000
rect 9404 132880 9456 132932
rect 9864 132880 9916 132932
rect 9128 132812 9180 132864
rect 319444 130364 319496 130416
rect 482652 130364 482704 130416
rect 5356 129820 5408 129872
rect 8208 129820 8260 129872
rect 356796 128596 356848 128648
rect 4528 127551 4580 127560
rect 4528 127517 4537 127551
rect 4537 127517 4571 127551
rect 4571 127517 4580 127551
rect 4528 127508 4580 127517
rect 5080 127372 5132 127424
rect 363604 126420 363656 126472
rect 312268 126284 312320 126336
rect 426624 126284 426676 126336
rect 477776 126123 477828 126132
rect 477776 126089 477785 126123
rect 477785 126089 477819 126123
rect 477819 126089 477828 126123
rect 477776 126080 477828 126089
rect 311532 125944 311584 125996
rect 312176 125944 312228 125996
rect 477684 125987 477736 125996
rect 477684 125953 477693 125987
rect 477693 125953 477727 125987
rect 477727 125953 477736 125987
rect 477684 125944 477736 125953
rect 3976 125536 4028 125588
rect 5356 125536 5408 125588
rect 428924 124899 428976 124908
rect 428924 124865 428933 124899
rect 428933 124865 428967 124899
rect 428967 124865 428976 124899
rect 428924 124856 428976 124865
rect 429200 124899 429252 124908
rect 429200 124865 429209 124899
rect 429209 124865 429243 124899
rect 429243 124865 429252 124899
rect 429200 124856 429252 124865
rect 429292 124899 429344 124908
rect 429292 124865 429301 124899
rect 429301 124865 429335 124899
rect 429335 124865 429344 124899
rect 429292 124856 429344 124865
rect 384304 124720 384356 124772
rect 360844 124652 360896 124704
rect 331864 123564 331916 123616
rect 366824 123403 366876 123412
rect 366824 123369 366833 123403
rect 366833 123369 366867 123403
rect 366867 123369 366876 123403
rect 366824 123360 366876 123369
rect 366732 123267 366784 123276
rect 366732 123233 366741 123267
rect 366741 123233 366775 123267
rect 366775 123233 366784 123267
rect 366732 123224 366784 123233
rect 367008 123199 367060 123208
rect 367008 123165 367017 123199
rect 367017 123165 367051 123199
rect 367051 123165 367060 123199
rect 367008 123156 367060 123165
rect 367100 123199 367152 123208
rect 367100 123165 367109 123199
rect 367109 123165 367143 123199
rect 367143 123165 367152 123199
rect 367100 123156 367152 123165
rect 318156 123020 318208 123072
rect 9128 121864 9180 121916
rect 385592 121864 385644 121916
rect 4068 121796 4120 121848
rect 321652 121796 321704 121848
rect 9496 121728 9548 121780
rect 311808 121728 311860 121780
rect 2780 121116 2832 121168
rect 5264 121116 5316 121168
rect 311992 120844 312044 120896
rect 7196 120776 7248 120828
rect 311072 120776 311124 120828
rect 20720 120708 20772 120760
rect 7104 120572 7156 120624
rect 129004 120708 129056 120760
rect 216128 120708 216180 120760
rect 310612 120708 310664 120760
rect 248880 120683 248932 120692
rect 248880 120649 248889 120683
rect 248889 120649 248923 120683
rect 248923 120649 248932 120683
rect 248880 120640 248932 120649
rect 299664 120683 299716 120692
rect 299664 120649 299673 120683
rect 299673 120649 299707 120683
rect 299707 120649 299716 120683
rect 299664 120640 299716 120649
rect 7012 120096 7064 120148
rect 221832 120096 221884 120148
rect 412088 120028 412140 120080
rect 5724 119960 5776 120012
rect 477684 119960 477736 120012
rect 451556 119892 451608 119944
rect 311164 119824 311216 119876
rect 311348 119688 311400 119740
rect 342076 119688 342128 119740
rect 216588 119620 216640 119672
rect 253940 119620 253992 119672
rect 254492 119620 254544 119672
rect 34980 119459 35032 119468
rect 34980 119425 34989 119459
rect 34989 119425 35023 119459
rect 35023 119425 35032 119459
rect 34980 119416 35032 119425
rect 35164 119459 35216 119468
rect 35164 119425 35173 119459
rect 35173 119425 35207 119459
rect 35207 119425 35216 119459
rect 35164 119416 35216 119425
rect 35348 119459 35400 119468
rect 35348 119425 35358 119459
rect 35358 119425 35392 119459
rect 35392 119425 35400 119459
rect 35348 119416 35400 119425
rect 38752 119459 38804 119468
rect 38752 119425 38761 119459
rect 38761 119425 38795 119459
rect 38795 119425 38804 119459
rect 38752 119416 38804 119425
rect 239128 119552 239180 119604
rect 239312 119552 239364 119604
rect 290556 119552 290608 119604
rect 290740 119552 290792 119604
rect 307668 119552 307720 119604
rect 308312 119620 308364 119672
rect 314200 119620 314252 119672
rect 310428 119552 310480 119604
rect 63500 119484 63552 119536
rect 63684 119459 63736 119468
rect 63684 119425 63693 119459
rect 63693 119425 63727 119459
rect 63727 119425 63736 119459
rect 63684 119416 63736 119425
rect 64052 119459 64104 119468
rect 64052 119425 64061 119459
rect 64061 119425 64095 119459
rect 64095 119425 64104 119459
rect 64052 119416 64104 119425
rect 145656 119459 145708 119468
rect 145656 119425 145665 119459
rect 145665 119425 145699 119459
rect 145699 119425 145708 119459
rect 145656 119416 145708 119425
rect 215576 119459 215628 119468
rect 162400 119391 162452 119400
rect 162400 119357 162409 119391
rect 162409 119357 162443 119391
rect 162443 119357 162452 119391
rect 162400 119348 162452 119357
rect 215576 119425 215585 119459
rect 215585 119425 215619 119459
rect 215619 119425 215628 119459
rect 215576 119416 215628 119425
rect 215760 119459 215812 119468
rect 215760 119425 215769 119459
rect 215769 119425 215803 119459
rect 215803 119425 215812 119459
rect 215760 119416 215812 119425
rect 215852 119459 215904 119468
rect 215852 119425 215861 119459
rect 215861 119425 215895 119459
rect 215895 119425 215904 119459
rect 216128 119459 216180 119468
rect 215852 119416 215904 119425
rect 216128 119425 216137 119459
rect 216137 119425 216171 119459
rect 216171 119425 216180 119459
rect 216128 119416 216180 119425
rect 216036 119391 216088 119400
rect 145748 119323 145800 119332
rect 145748 119289 145757 119323
rect 145757 119289 145791 119323
rect 145791 119289 145800 119323
rect 145748 119280 145800 119289
rect 216036 119357 216045 119391
rect 216045 119357 216079 119391
rect 216079 119357 216088 119391
rect 216036 119348 216088 119357
rect 238760 119459 238812 119468
rect 238760 119425 238769 119459
rect 238769 119425 238803 119459
rect 238803 119425 238812 119459
rect 238760 119416 238812 119425
rect 238852 119459 238904 119468
rect 238852 119425 238861 119459
rect 238861 119425 238895 119459
rect 238895 119425 238904 119459
rect 239404 119484 239456 119536
rect 289912 119484 289964 119536
rect 254216 119459 254268 119468
rect 238852 119416 238904 119425
rect 254216 119425 254225 119459
rect 254225 119425 254259 119459
rect 254259 119425 254268 119459
rect 254216 119416 254268 119425
rect 289728 119416 289780 119468
rect 290464 119484 290516 119536
rect 5908 119212 5960 119264
rect 34888 119255 34940 119264
rect 34888 119221 34897 119255
rect 34897 119221 34931 119255
rect 34931 119221 34940 119255
rect 34888 119212 34940 119221
rect 38844 119255 38896 119264
rect 38844 119221 38853 119255
rect 38853 119221 38887 119255
rect 38887 119221 38896 119255
rect 38844 119212 38896 119221
rect 161020 119255 161072 119264
rect 161020 119221 161029 119255
rect 161029 119221 161063 119255
rect 161063 119221 161072 119255
rect 161020 119212 161072 119221
rect 172704 119255 172756 119264
rect 172704 119221 172713 119255
rect 172713 119221 172747 119255
rect 172747 119221 172756 119255
rect 172704 119212 172756 119221
rect 239036 119348 239088 119400
rect 239312 119348 239364 119400
rect 248512 119348 248564 119400
rect 238944 119212 238996 119264
rect 248236 119212 248288 119264
rect 290372 119348 290424 119400
rect 434720 119484 434772 119536
rect 292120 119348 292172 119400
rect 385776 119416 385828 119468
rect 355508 119348 355560 119400
rect 351920 119280 351972 119332
rect 496544 119212 496596 119264
rect 34612 119051 34664 119060
rect 34612 119017 34621 119051
rect 34621 119017 34655 119051
rect 34655 119017 34664 119051
rect 34612 119008 34664 119017
rect 48136 119008 48188 119060
rect 4896 118940 4948 118992
rect 145656 118940 145708 118992
rect 157524 118940 157576 118992
rect 168104 118940 168156 118992
rect 238760 119008 238812 119060
rect 290740 119076 290792 119128
rect 340972 119144 341024 119196
rect 313740 119076 313792 119128
rect 318156 119008 318208 119060
rect 179328 118872 179380 118924
rect 34796 118847 34848 118856
rect 34796 118813 34805 118847
rect 34805 118813 34839 118847
rect 34839 118813 34848 118847
rect 34796 118804 34848 118813
rect 34888 118847 34940 118856
rect 34888 118813 34897 118847
rect 34897 118813 34931 118847
rect 34931 118813 34940 118847
rect 35164 118847 35216 118856
rect 34888 118804 34940 118813
rect 35164 118813 35173 118847
rect 35173 118813 35207 118847
rect 35207 118813 35216 118847
rect 35164 118804 35216 118813
rect 162400 118804 162452 118856
rect 180892 118804 180944 118856
rect 238852 118872 238904 118924
rect 317972 118940 318024 118992
rect 318616 118804 318668 118856
rect 311624 118736 311676 118788
rect 317696 118668 317748 118720
rect 9680 118600 9732 118652
rect 23020 118600 23072 118652
rect 56232 118600 56284 118652
rect 496268 118600 496320 118652
rect 4620 118532 4672 118584
rect 16764 118532 16816 118584
rect 155592 118532 155644 118584
rect 496176 118532 496228 118584
rect 162216 118464 162268 118516
rect 496636 118464 496688 118516
rect 3700 118396 3752 118448
rect 4896 118396 4948 118448
rect 282000 118396 282052 118448
rect 467840 118396 467892 118448
rect 202236 118328 202288 118380
rect 496084 118328 496136 118380
rect 6276 118260 6328 118312
rect 215484 118260 215536 118312
rect 222108 118260 222160 118312
rect 444012 118260 444064 118312
rect 228824 118192 228876 118244
rect 438308 118192 438360 118244
rect 209136 118124 209188 118176
rect 412640 118124 412692 118176
rect 122196 118056 122248 118108
rect 122748 118056 122800 118108
rect 316776 118056 316828 118108
rect 308496 117988 308548 118040
rect 409420 117988 409472 118040
rect 10416 117920 10468 117972
rect 384304 117920 384356 117972
rect 175924 117852 175976 117904
rect 316868 117852 316920 117904
rect 195336 117784 195388 117836
rect 316960 117784 317012 117836
rect 295156 117716 295208 117768
rect 369860 117716 369912 117768
rect 6184 117648 6236 117700
rect 301596 117648 301648 117700
rect 310980 117648 311032 117700
rect 70032 117580 70084 117632
rect 310428 117580 310480 117632
rect 22100 117308 22152 117360
rect 23020 117308 23072 117360
rect 89260 117308 89312 117360
rect 106464 117308 106516 117360
rect 451372 117283 451424 117292
rect 451372 117249 451390 117283
rect 451390 117249 451424 117283
rect 451372 117240 451424 117249
rect 451648 117283 451700 117292
rect 451648 117249 451657 117283
rect 451657 117249 451691 117283
rect 451691 117249 451700 117283
rect 451648 117240 451700 117249
rect 314108 117036 314160 117088
rect 450268 117079 450320 117088
rect 450268 117045 450277 117079
rect 450277 117045 450311 117079
rect 450311 117045 450320 117079
rect 450268 117036 450320 117045
rect 314568 116628 314620 116680
rect 209504 116560 209556 116612
rect 310796 116560 310848 116612
rect 451648 116560 451700 116612
rect 458180 116560 458232 116612
rect 495440 116560 495492 116612
rect 209504 115787 209556 115796
rect 209504 115753 209513 115787
rect 209513 115753 209547 115787
rect 209547 115753 209556 115787
rect 209504 115744 209556 115753
rect 209872 115651 209924 115660
rect 209872 115617 209881 115651
rect 209881 115617 209915 115651
rect 209915 115617 209924 115651
rect 209872 115608 209924 115617
rect 209688 115583 209740 115592
rect 209688 115549 209697 115583
rect 209697 115549 209731 115583
rect 209731 115549 209740 115583
rect 209688 115540 209740 115549
rect 328552 115540 328604 115592
rect 315396 114860 315448 114912
rect 89260 113976 89312 114028
rect 32496 113883 32548 113892
rect 32496 113849 32505 113883
rect 32505 113849 32539 113883
rect 32539 113849 32548 113883
rect 32496 113840 32548 113849
rect 69388 113407 69440 113416
rect 69388 113373 69397 113407
rect 69397 113373 69431 113407
rect 69431 113373 69440 113407
rect 69388 113364 69440 113373
rect 310244 113364 310296 113416
rect 346768 113228 346820 113280
rect 273260 112956 273312 113008
rect 405740 112956 405792 113008
rect 260288 112888 260340 112940
rect 460204 112888 460256 112940
rect 266912 112820 266964 112872
rect 405832 112820 405884 112872
rect 121184 112752 121236 112804
rect 396724 112752 396776 112804
rect 127808 112684 127860 112736
rect 418712 112684 418764 112736
rect 28448 112548 28500 112600
rect 319444 112548 319496 112600
rect 81440 112480 81492 112532
rect 403348 112480 403400 112532
rect 48320 112412 48372 112464
rect 380164 112412 380216 112464
rect 15200 112344 15252 112396
rect 370504 112344 370556 112396
rect 316684 112276 316736 112328
rect 327356 112276 327408 112328
rect 328552 112251 328604 112260
rect 293408 112140 293460 112192
rect 328276 112183 328328 112192
rect 220544 111936 220596 111988
rect 327908 112004 327960 112056
rect 328276 112149 328285 112183
rect 328285 112149 328319 112183
rect 328319 112149 328328 112183
rect 328276 112140 328328 112149
rect 328552 112217 328561 112251
rect 328561 112217 328595 112251
rect 328595 112217 328604 112251
rect 328552 112208 328604 112217
rect 489920 112140 489972 112192
rect 456064 111936 456116 111988
rect 114560 111868 114612 111920
rect 115112 111868 115164 111920
rect 393320 111868 393372 111920
rect 327264 111843 327316 111852
rect 327264 111809 327273 111843
rect 327273 111809 327307 111843
rect 327307 111809 327316 111843
rect 327264 111800 327316 111809
rect 327356 111843 327408 111852
rect 327356 111809 327365 111843
rect 327365 111809 327399 111843
rect 327399 111809 327408 111843
rect 328552 111843 328604 111852
rect 327356 111800 327408 111809
rect 328552 111809 328561 111843
rect 328561 111809 328595 111843
rect 328595 111809 328604 111843
rect 328552 111800 328604 111809
rect 337476 111800 337528 111852
rect 494060 111732 494112 111784
rect 183468 111664 183520 111716
rect 419632 111664 419684 111716
rect 168104 111596 168156 111648
rect 194508 111596 194560 111648
rect 9036 111528 9088 111580
rect 132776 111528 132828 111580
rect 135720 111528 135772 111580
rect 214564 111528 214616 111580
rect 341432 111596 341484 111648
rect 480628 111639 480680 111648
rect 480628 111605 480637 111639
rect 480637 111605 480671 111639
rect 480671 111605 480680 111639
rect 480628 111596 480680 111605
rect 209688 111392 209740 111444
rect 416412 111392 416464 111444
rect 5632 111324 5684 111376
rect 181352 111324 181404 111376
rect 106464 111256 106516 111308
rect 162400 111256 162452 111308
rect 168380 111256 168432 111308
rect 181628 111256 181680 111308
rect 222384 111324 222436 111376
rect 417424 111324 417476 111376
rect 6644 111188 6696 111240
rect 181812 111120 181864 111172
rect 182088 111188 182140 111240
rect 182824 111188 182876 111240
rect 367100 111256 367152 111308
rect 213644 111188 213696 111240
rect 221924 111188 221976 111240
rect 222016 111188 222068 111240
rect 231860 111120 231912 111172
rect 310336 111120 310388 111172
rect 472624 111188 472676 111240
rect 179328 111095 179380 111104
rect 179328 111061 179337 111095
rect 179337 111061 179371 111095
rect 179371 111061 179380 111095
rect 179328 111052 179380 111061
rect 179880 111052 179932 111104
rect 316592 111052 316644 111104
rect 183192 110984 183244 111036
rect 183100 110916 183152 110968
rect 202512 110848 202564 110900
rect 203064 110848 203116 110900
rect 5264 110780 5316 110832
rect 274180 110984 274232 111036
rect 273444 110848 273496 110900
rect 274640 110848 274692 110900
rect 314108 110984 314160 111036
rect 315396 110916 315448 110968
rect 495440 110780 495492 110832
rect 96896 110755 96948 110764
rect 35164 110644 35216 110696
rect 96896 110721 96905 110755
rect 96905 110721 96939 110755
rect 96939 110721 96948 110755
rect 96896 110712 96948 110721
rect 106464 110755 106516 110764
rect 106464 110721 106473 110755
rect 106473 110721 106507 110755
rect 106507 110721 106516 110755
rect 106464 110712 106516 110721
rect 168104 110755 168156 110764
rect 168104 110721 168113 110755
rect 168113 110721 168147 110755
rect 168147 110721 168156 110755
rect 168104 110712 168156 110721
rect 168380 110712 168432 110764
rect 180616 110755 180668 110764
rect 180616 110721 180634 110755
rect 180634 110721 180668 110755
rect 182640 110755 182692 110764
rect 180616 110712 180668 110721
rect 182640 110721 182649 110755
rect 182649 110721 182683 110755
rect 182683 110721 182692 110755
rect 182640 110712 182692 110721
rect 194324 110712 194376 110764
rect 194416 110755 194468 110764
rect 194416 110721 194425 110755
rect 194425 110721 194459 110755
rect 194459 110721 194468 110755
rect 194416 110712 194468 110721
rect 194600 110712 194652 110764
rect 194692 110712 194744 110764
rect 214380 110712 214432 110764
rect 214472 110755 214524 110764
rect 214472 110721 214481 110755
rect 214481 110721 214515 110755
rect 214515 110721 214524 110755
rect 214656 110755 214708 110764
rect 214472 110712 214524 110721
rect 214656 110721 214665 110755
rect 214665 110721 214699 110755
rect 214699 110721 214708 110755
rect 214656 110712 214708 110721
rect 222016 110755 222068 110764
rect 222016 110721 222024 110755
rect 222024 110721 222058 110755
rect 222058 110721 222068 110755
rect 222016 110712 222068 110721
rect 222200 110755 222252 110764
rect 222200 110721 222209 110755
rect 222209 110721 222243 110755
rect 222243 110721 222252 110755
rect 222200 110712 222252 110721
rect 222384 110755 222436 110764
rect 222384 110721 222393 110755
rect 222393 110721 222427 110755
rect 222427 110721 222436 110755
rect 222384 110712 222436 110721
rect 222568 110712 222620 110764
rect 418988 110712 419040 110764
rect 179880 110644 179932 110696
rect 180892 110687 180944 110696
rect 180892 110653 180901 110687
rect 180901 110653 180935 110687
rect 180935 110653 180944 110687
rect 180892 110644 180944 110653
rect 181260 110644 181312 110696
rect 182088 110687 182140 110696
rect 182088 110653 182097 110687
rect 182097 110653 182131 110687
rect 182131 110653 182140 110687
rect 182088 110644 182140 110653
rect 222108 110687 222160 110696
rect 222108 110653 222112 110687
rect 222112 110653 222146 110687
rect 222146 110653 222160 110687
rect 222108 110644 222160 110653
rect 6828 110576 6880 110628
rect 4988 110508 5040 110560
rect 168104 110619 168156 110628
rect 137192 110551 137244 110560
rect 137192 110517 137201 110551
rect 137201 110517 137235 110551
rect 137235 110517 137244 110551
rect 137192 110508 137244 110517
rect 168104 110585 168113 110619
rect 168113 110585 168147 110619
rect 168147 110585 168156 110619
rect 168104 110576 168156 110585
rect 170220 110551 170272 110560
rect 170220 110517 170229 110551
rect 170229 110517 170263 110551
rect 170263 110517 170272 110551
rect 170220 110508 170272 110517
rect 179512 110551 179564 110560
rect 179512 110517 179521 110551
rect 179521 110517 179555 110551
rect 179555 110517 179564 110551
rect 179512 110508 179564 110517
rect 190460 110551 190512 110560
rect 190460 110517 190469 110551
rect 190469 110517 190503 110551
rect 190503 110517 190512 110551
rect 190460 110508 190512 110517
rect 273444 110644 273496 110696
rect 273628 110687 273680 110696
rect 273628 110653 273637 110687
rect 273637 110653 273671 110687
rect 273671 110653 273680 110687
rect 273628 110644 273680 110653
rect 273812 110687 273864 110696
rect 273812 110653 273821 110687
rect 273821 110653 273855 110687
rect 273855 110653 273864 110687
rect 273812 110644 273864 110653
rect 409052 110644 409104 110696
rect 214380 110551 214432 110560
rect 214380 110517 214389 110551
rect 214389 110517 214423 110551
rect 214423 110517 214432 110551
rect 214380 110508 214432 110517
rect 214472 110508 214524 110560
rect 222384 110508 222436 110560
rect 310888 110576 310940 110628
rect 273168 110551 273220 110560
rect 273168 110517 273177 110551
rect 273177 110517 273211 110551
rect 273211 110517 273220 110551
rect 273168 110508 273220 110517
rect 311164 110508 311216 110560
rect 273444 110304 273496 110356
rect 8576 109692 8628 109744
rect 22100 109692 22152 109744
rect 8484 109284 8536 109336
rect 20720 109284 20772 109336
rect 21548 109284 21600 109336
rect 7012 109148 7064 109200
rect 8668 109148 8720 109200
rect 8668 109012 8720 109064
rect 180892 109284 180944 109336
rect 453028 109191 453080 109200
rect 453028 109157 453037 109191
rect 453037 109157 453071 109191
rect 453071 109157 453080 109191
rect 453028 109148 453080 109157
rect 470600 109012 470652 109064
rect 5080 108536 5132 108588
rect 315212 108536 315264 108588
rect 8944 108468 8996 108520
rect 366732 108468 366784 108520
rect 8392 108400 8444 108452
rect 368020 108400 368072 108452
rect 7104 108332 7156 108384
rect 491300 108332 491352 108384
rect 5172 108264 5224 108316
rect 416596 108264 416648 108316
rect 317236 107924 317288 107976
rect 419540 107967 419592 107976
rect 419540 107933 419549 107967
rect 419549 107933 419583 107967
rect 419583 107933 419592 107967
rect 419540 107924 419592 107933
rect 471888 107924 471940 107976
rect 317052 107788 317104 107840
rect 9496 107652 9548 107704
rect 312728 107652 312780 107704
rect 358084 106292 358136 106344
rect 368388 105451 368440 105460
rect 368388 105417 368397 105451
rect 368397 105417 368431 105451
rect 368431 105417 368440 105451
rect 368388 105408 368440 105417
rect 372620 105272 372672 105324
rect 317972 105068 318024 105120
rect 368388 105068 368440 105120
rect 344652 102144 344704 102196
rect 495532 102144 495584 102196
rect 2964 101056 3016 101108
rect 3700 101099 3752 101108
rect 3700 101065 3709 101099
rect 3709 101065 3743 101099
rect 3743 101065 3752 101099
rect 3700 101056 3752 101065
rect 9496 100988 9548 101040
rect 4988 100784 5040 100836
rect 3332 100759 3384 100768
rect 3332 100725 3341 100759
rect 3341 100725 3375 100759
rect 3375 100725 3384 100759
rect 3332 100716 3384 100725
rect 5264 100716 5316 100768
rect 6184 100716 6236 100768
rect 388444 100716 388496 100768
rect 396632 99220 396684 99272
rect 458180 99263 458232 99272
rect 440884 99152 440936 99204
rect 458180 99229 458189 99263
rect 458189 99229 458223 99263
rect 458223 99229 458232 99263
rect 458180 99220 458232 99229
rect 495532 99220 495584 99272
rect 456800 99127 456852 99136
rect 456800 99093 456809 99127
rect 456809 99093 456843 99127
rect 456843 99093 456852 99127
rect 456800 99084 456852 99093
rect 432604 93780 432656 93832
rect 495532 93780 495584 93832
rect 436744 90108 436796 90160
rect 433984 90040 434036 90092
rect 318616 89836 318668 89888
rect 439964 89879 440016 89888
rect 439964 89845 439973 89879
rect 439973 89845 440007 89879
rect 440007 89845 440016 89879
rect 439964 89836 440016 89845
rect 5356 89632 5408 89684
rect 8024 89632 8076 89684
rect 348424 89632 348476 89684
rect 495532 89632 495584 89684
rect 312544 85756 312596 85808
rect 382188 85756 382240 85808
rect 312820 85688 312872 85740
rect 327724 85552 327776 85604
rect 311992 85484 312044 85536
rect 312912 85484 312964 85536
rect 318064 84736 318116 84788
rect 369124 84600 369176 84652
rect 8852 79883 8904 79892
rect 8852 79849 8861 79883
rect 8861 79849 8895 79883
rect 8895 79849 8904 79883
rect 8852 79840 8904 79849
rect 9128 79772 9180 79824
rect 6184 79704 6236 79756
rect 8944 79679 8996 79688
rect 8944 79645 8953 79679
rect 8953 79645 8987 79679
rect 8987 79645 8996 79679
rect 8944 79636 8996 79645
rect 9128 79679 9180 79688
rect 9128 79645 9137 79679
rect 9137 79645 9171 79679
rect 9171 79645 9180 79679
rect 9128 79636 9180 79645
rect 8300 79568 8352 79620
rect 443092 79271 443144 79280
rect 443092 79237 443101 79271
rect 443101 79237 443135 79271
rect 443135 79237 443144 79271
rect 443092 79228 443144 79237
rect 442908 79203 442960 79212
rect 442908 79169 442917 79203
rect 442917 79169 442951 79203
rect 442951 79169 442960 79203
rect 442908 79160 442960 79169
rect 443184 78999 443236 79008
rect 443184 78965 443193 78999
rect 443193 78965 443227 78999
rect 443227 78965 443236 78999
rect 443184 78956 443236 78965
rect 337752 78659 337804 78668
rect 337752 78625 337761 78659
rect 337761 78625 337795 78659
rect 337795 78625 337804 78659
rect 338212 78659 338264 78668
rect 337752 78616 337804 78625
rect 338212 78625 338221 78659
rect 338221 78625 338255 78659
rect 338255 78625 338264 78659
rect 338212 78616 338264 78625
rect 429844 78616 429896 78668
rect 469864 78659 469916 78668
rect 469864 78625 469873 78659
rect 469873 78625 469907 78659
rect 469907 78625 469916 78659
rect 469864 78616 469916 78625
rect 327816 78548 327868 78600
rect 338028 78591 338080 78600
rect 338028 78557 338037 78591
rect 338037 78557 338071 78591
rect 338071 78557 338080 78591
rect 338028 78548 338080 78557
rect 339316 78548 339368 78600
rect 469588 78591 469640 78600
rect 469588 78557 469597 78591
rect 469597 78557 469631 78591
rect 469631 78557 469640 78591
rect 469588 78548 469640 78557
rect 469680 78591 469732 78600
rect 469680 78557 469689 78591
rect 469689 78557 469723 78591
rect 469723 78557 469732 78591
rect 469680 78548 469732 78557
rect 473728 78548 473780 78600
rect 406384 78480 406436 78532
rect 469404 78455 469456 78464
rect 469404 78421 469413 78455
rect 469413 78421 469447 78455
rect 469447 78421 469456 78455
rect 469404 78412 469456 78421
rect 442540 78208 442592 78260
rect 2780 76916 2832 76968
rect 4712 76916 4764 76968
rect 429844 75531 429896 75540
rect 429844 75497 429853 75531
rect 429853 75497 429887 75531
rect 429887 75497 429896 75531
rect 429844 75488 429896 75497
rect 429660 75327 429712 75336
rect 429660 75293 429669 75327
rect 429669 75293 429703 75327
rect 429703 75293 429712 75327
rect 429660 75284 429712 75293
rect 362224 72632 362276 72684
rect 370504 72564 370556 72616
rect 378968 72607 379020 72616
rect 378968 72573 378977 72607
rect 378977 72573 379011 72607
rect 379011 72573 379020 72607
rect 378968 72564 379020 72573
rect 367468 72428 367520 72480
rect 378968 72428 379020 72480
rect 382188 72428 382240 72480
rect 418436 72428 418488 72480
rect 496452 72267 496504 72276
rect 496452 72233 496461 72267
rect 496461 72233 496495 72267
rect 496495 72233 496504 72267
rect 496452 72224 496504 72233
rect 359464 70388 359516 70440
rect 376208 67532 376260 67584
rect 376668 67532 376720 67584
rect 429660 67532 429712 67584
rect 310060 67371 310112 67380
rect 310060 67337 310069 67371
rect 310069 67337 310103 67371
rect 310103 67337 310112 67371
rect 310060 67328 310112 67337
rect 339316 67192 339368 67244
rect 314108 66580 314160 66632
rect 376668 66580 376720 66632
rect 360108 66487 360160 66496
rect 360108 66453 360117 66487
rect 360117 66453 360151 66487
rect 360151 66453 360160 66487
rect 360108 66444 360160 66453
rect 445760 66444 445812 66496
rect 9220 66104 9272 66156
rect 9036 65968 9088 66020
rect 493876 65535 493928 65544
rect 493876 65501 493885 65535
rect 493885 65501 493919 65535
rect 493919 65501 493928 65535
rect 493876 65492 493928 65501
rect 314016 63724 314068 63776
rect 480628 63452 480680 63504
rect 495532 63452 495584 63504
rect 344928 61208 344980 61260
rect 446036 61251 446088 61260
rect 446036 61217 446045 61251
rect 446045 61217 446079 61251
rect 446079 61217 446088 61251
rect 446036 61208 446088 61217
rect 445668 61183 445720 61192
rect 445668 61149 445677 61183
rect 445677 61149 445711 61183
rect 445711 61149 445720 61183
rect 445668 61140 445720 61149
rect 445760 61183 445812 61192
rect 445760 61149 445769 61183
rect 445769 61149 445803 61183
rect 445803 61149 445812 61183
rect 445760 61140 445812 61149
rect 496084 61072 496136 61124
rect 422944 61004 422996 61056
rect 406292 59712 406344 59764
rect 443184 59712 443236 59764
rect 315396 59576 315448 59628
rect 419540 59644 419592 59696
rect 372712 59619 372764 59628
rect 372712 59585 372721 59619
rect 372721 59585 372755 59619
rect 372755 59585 372764 59619
rect 372712 59576 372764 59585
rect 406292 59619 406344 59628
rect 406292 59585 406301 59619
rect 406301 59585 406335 59619
rect 406335 59585 406344 59619
rect 406292 59576 406344 59585
rect 401232 59508 401284 59560
rect 406476 59619 406528 59628
rect 406476 59585 406486 59619
rect 406486 59585 406520 59619
rect 406520 59585 406528 59619
rect 406476 59576 406528 59585
rect 464252 59576 464304 59628
rect 344284 59440 344336 59492
rect 342904 59372 342956 59424
rect 398104 59168 398156 59220
rect 495532 59168 495584 59220
rect 7104 58488 7156 58540
rect 2780 58216 2832 58268
rect 5172 58216 5224 58268
rect 313740 57400 313792 57452
rect 318156 57196 318208 57248
rect 422024 57239 422076 57248
rect 422024 57205 422033 57239
rect 422033 57205 422067 57239
rect 422067 57205 422076 57239
rect 422024 57196 422076 57205
rect 312452 55836 312504 55888
rect 320180 55836 320232 55888
rect 9404 54816 9456 54868
rect 401232 54655 401284 54664
rect 401232 54621 401241 54655
rect 401241 54621 401275 54655
rect 401275 54621 401284 54655
rect 401232 54612 401284 54621
rect 401140 54519 401192 54528
rect 401140 54485 401149 54519
rect 401149 54485 401183 54519
rect 401183 54485 401192 54519
rect 401140 54476 401192 54485
rect 442908 54476 442960 54528
rect 2780 53660 2832 53712
rect 5080 53660 5132 53712
rect 367008 50260 367060 50312
rect 385224 50124 385276 50176
rect 311716 48220 311768 48272
rect 463884 48127 463936 48136
rect 463884 48093 463893 48127
rect 463893 48093 463927 48127
rect 463927 48093 463936 48127
rect 463884 48084 463936 48093
rect 314476 46316 314528 46368
rect 318524 46044 318576 46096
rect 318708 45976 318760 46028
rect 430580 45976 430632 46028
rect 339960 45951 340012 45960
rect 339960 45917 339969 45951
rect 339969 45917 340003 45951
rect 340003 45917 340012 45951
rect 339960 45908 340012 45917
rect 318064 45772 318116 45824
rect 340420 45772 340472 45824
rect 369216 45500 369268 45552
rect 495532 45500 495584 45552
rect 311900 45024 311952 45076
rect 310152 44888 310204 44940
rect 378968 44888 379020 44940
rect 310428 44863 310480 44872
rect 310428 44829 310437 44863
rect 310437 44829 310471 44863
rect 310471 44829 310480 44863
rect 310428 44820 310480 44829
rect 310244 44684 310296 44736
rect 496360 43052 496412 43104
rect 8392 42236 8444 42288
rect 8024 42143 8076 42152
rect 8024 42109 8033 42143
rect 8033 42109 8067 42143
rect 8067 42109 8076 42143
rect 8024 42100 8076 42109
rect 9404 42007 9456 42016
rect 9404 41973 9413 42007
rect 9413 41973 9447 42007
rect 9447 41973 9456 42007
rect 9404 41964 9456 41973
rect 338764 39788 338816 39840
rect 384304 37816 384356 37868
rect 418344 37791 418396 37800
rect 418344 37757 418353 37791
rect 418353 37757 418387 37791
rect 418387 37757 418396 37791
rect 418344 37748 418396 37757
rect 418436 37791 418488 37800
rect 418436 37757 418445 37791
rect 418445 37757 418479 37791
rect 418479 37757 418488 37791
rect 418436 37748 418488 37757
rect 479432 37748 479484 37800
rect 395344 37612 395396 37664
rect 417884 37655 417936 37664
rect 417884 37621 417893 37655
rect 417893 37621 417927 37655
rect 417927 37621 417936 37655
rect 417884 37612 417936 37621
rect 312728 36660 312780 36712
rect 368480 36660 368532 36712
rect 312636 36592 312688 36644
rect 463884 36592 463936 36644
rect 311624 36524 311676 36576
rect 466460 36524 466512 36576
rect 346492 36320 346544 36372
rect 343916 36159 343968 36168
rect 343916 36125 343925 36159
rect 343925 36125 343959 36159
rect 343959 36125 343968 36159
rect 343916 36116 343968 36125
rect 373172 36116 373224 36168
rect 346308 36048 346360 36100
rect 410524 35844 410576 35896
rect 495532 35844 495584 35896
rect 390928 35275 390980 35284
rect 390928 35241 390937 35275
rect 390937 35241 390971 35275
rect 390971 35241 390980 35275
rect 390928 35232 390980 35241
rect 392032 35071 392084 35080
rect 392032 35037 392050 35071
rect 392050 35037 392084 35071
rect 392032 35028 392084 35037
rect 416872 35028 416924 35080
rect 371792 34731 371844 34740
rect 371792 34697 371801 34731
rect 371801 34697 371835 34731
rect 371835 34697 371844 34731
rect 371792 34688 371844 34697
rect 372896 34595 372948 34604
rect 372896 34561 372914 34595
rect 372914 34561 372948 34595
rect 372896 34552 372948 34561
rect 373172 34595 373224 34604
rect 373172 34561 373181 34595
rect 373181 34561 373215 34595
rect 373215 34561 373224 34595
rect 373172 34552 373224 34561
rect 399484 32011 399536 32020
rect 399484 31977 399493 32011
rect 399493 31977 399527 32011
rect 399527 31977 399536 32011
rect 399484 31968 399536 31977
rect 321376 31424 321428 31476
rect 416688 31424 416740 31476
rect 417516 31467 417568 31476
rect 417516 31433 417525 31467
rect 417525 31433 417559 31467
rect 417559 31433 417568 31467
rect 417516 31424 417568 31433
rect 416872 31356 416924 31408
rect 416872 31263 416924 31272
rect 416872 31229 416881 31263
rect 416881 31229 416915 31263
rect 416915 31229 416924 31263
rect 416872 31220 416924 31229
rect 458180 31220 458232 31272
rect 415492 31127 415544 31136
rect 415492 31093 415501 31127
rect 415501 31093 415535 31127
rect 415535 31093 415544 31127
rect 415492 31084 415544 31093
rect 463516 31084 463568 31136
rect 311348 30676 311400 30728
rect 318340 30268 318392 30320
rect 320456 30311 320508 30320
rect 320456 30277 320465 30311
rect 320465 30277 320499 30311
rect 320499 30277 320508 30311
rect 320456 30268 320508 30277
rect 318432 30200 318484 30252
rect 376024 27455 376076 27464
rect 376024 27421 376033 27455
rect 376033 27421 376067 27455
rect 376067 27421 376076 27455
rect 376024 27412 376076 27421
rect 9312 25891 9364 25900
rect 9312 25857 9321 25891
rect 9321 25857 9355 25891
rect 9355 25857 9364 25891
rect 9312 25848 9364 25857
rect 9496 25823 9548 25832
rect 9496 25789 9505 25823
rect 9505 25789 9539 25823
rect 9539 25789 9548 25823
rect 9496 25780 9548 25789
rect 9220 25644 9272 25696
rect 310152 25347 310204 25356
rect 310152 25313 310161 25347
rect 310161 25313 310195 25347
rect 310195 25313 310204 25347
rect 310152 25304 310204 25313
rect 310612 25304 310664 25356
rect 311532 25236 311584 25288
rect 360200 25100 360252 25152
rect 356704 23400 356756 23452
rect 495532 23400 495584 23452
rect 456064 16099 456116 16108
rect 456064 16065 456073 16099
rect 456073 16065 456107 16099
rect 456107 16065 456116 16099
rect 456064 16056 456116 16065
rect 317144 15852 317196 15904
rect 318248 15444 318300 15496
rect 315672 15376 315724 15428
rect 453028 15444 453080 15496
rect 496360 15487 496412 15496
rect 496360 15453 496369 15487
rect 496369 15453 496403 15487
rect 496403 15453 496412 15487
rect 496360 15444 496412 15453
rect 335544 15308 335596 15360
rect 335636 15308 335688 15360
rect 447784 15308 447836 15360
rect 475384 14016 475436 14068
rect 460204 13948 460256 14000
rect 414664 13812 414716 13864
rect 479432 13855 479484 13864
rect 479432 13821 479441 13855
rect 479441 13821 479475 13855
rect 479475 13821 479484 13855
rect 479432 13812 479484 13821
rect 351184 13744 351236 13796
rect 495440 13744 495492 13796
rect 344652 12427 344704 12436
rect 344652 12393 344661 12427
rect 344661 12393 344695 12427
rect 344695 12393 344704 12427
rect 344652 12384 344704 12393
rect 9496 11840 9548 11892
rect 417884 11840 417936 11892
rect 261852 10616 261904 10668
rect 315488 10616 315540 10668
rect 239956 10548 240008 10600
rect 310152 10548 310204 10600
rect 244648 10480 244700 10532
rect 450268 10480 450320 10532
rect 147956 10412 148008 10464
rect 371792 10412 371844 10464
rect 116768 10344 116820 10396
rect 342352 10344 342404 10396
rect 151268 10276 151320 10328
rect 383752 10276 383804 10328
rect 168656 9868 168708 9920
rect 169116 9868 169168 9920
rect 151268 9707 151320 9716
rect 77300 9596 77352 9648
rect 151268 9673 151277 9707
rect 151277 9673 151311 9707
rect 151311 9673 151320 9707
rect 151268 9664 151320 9673
rect 168656 9664 168708 9716
rect 8760 9528 8812 9580
rect 77116 9571 77168 9580
rect 77116 9537 77125 9571
rect 77125 9537 77159 9571
rect 77159 9537 77168 9571
rect 77116 9528 77168 9537
rect 77852 9571 77904 9580
rect 77852 9537 77861 9571
rect 77861 9537 77895 9571
rect 77895 9537 77904 9571
rect 77852 9528 77904 9537
rect 78588 9596 78640 9648
rect 168932 9664 168984 9716
rect 168840 9596 168892 9648
rect 169116 9634 169168 9686
rect 239956 9707 240008 9716
rect 239956 9673 239965 9707
rect 239965 9673 239999 9707
rect 239999 9673 240008 9707
rect 239956 9664 240008 9673
rect 248144 9707 248196 9716
rect 248144 9673 248153 9707
rect 248153 9673 248187 9707
rect 248187 9673 248196 9707
rect 248144 9664 248196 9673
rect 272340 9664 272392 9716
rect 277768 9707 277820 9716
rect 272156 9596 272208 9648
rect 78864 9571 78916 9580
rect 78864 9537 78873 9571
rect 78873 9537 78907 9571
rect 78907 9537 78916 9571
rect 78864 9528 78916 9537
rect 79048 9571 79100 9580
rect 79048 9537 79057 9571
rect 79057 9537 79091 9571
rect 79091 9537 79100 9571
rect 88432 9571 88484 9580
rect 79048 9528 79100 9537
rect 88432 9537 88441 9571
rect 88441 9537 88475 9571
rect 88475 9537 88484 9571
rect 88432 9528 88484 9537
rect 88616 9571 88668 9580
rect 88616 9537 88625 9571
rect 88625 9537 88659 9571
rect 88659 9537 88668 9571
rect 88616 9528 88668 9537
rect 95148 9571 95200 9580
rect 95148 9537 95157 9571
rect 95157 9537 95191 9571
rect 95191 9537 95200 9571
rect 95148 9528 95200 9537
rect 116492 9571 116544 9580
rect 79232 9503 79284 9512
rect 7748 9392 7800 9444
rect 65156 9435 65208 9444
rect 65156 9401 65165 9435
rect 65165 9401 65199 9435
rect 65199 9401 65208 9435
rect 65156 9392 65208 9401
rect 79232 9469 79241 9503
rect 79241 9469 79275 9503
rect 79275 9469 79284 9503
rect 79232 9460 79284 9469
rect 88340 9435 88392 9444
rect 2780 9324 2832 9376
rect 4804 9324 4856 9376
rect 35532 9367 35584 9376
rect 35532 9333 35541 9367
rect 35541 9333 35575 9367
rect 35575 9333 35584 9367
rect 35532 9324 35584 9333
rect 72240 9367 72292 9376
rect 72240 9333 72249 9367
rect 72249 9333 72283 9367
rect 72283 9333 72292 9367
rect 72240 9324 72292 9333
rect 77944 9367 77996 9376
rect 77944 9333 77953 9367
rect 77953 9333 77987 9367
rect 77987 9333 77996 9367
rect 77944 9324 77996 9333
rect 88340 9401 88349 9435
rect 88349 9401 88383 9435
rect 88383 9401 88392 9435
rect 88340 9392 88392 9401
rect 116492 9537 116501 9571
rect 116501 9537 116535 9571
rect 116535 9537 116544 9571
rect 116492 9528 116544 9537
rect 116584 9571 116636 9580
rect 116584 9537 116593 9571
rect 116593 9537 116627 9571
rect 116627 9537 116636 9571
rect 116768 9571 116820 9580
rect 116584 9528 116636 9537
rect 116768 9537 116777 9571
rect 116777 9537 116811 9571
rect 116811 9537 116820 9571
rect 116768 9528 116820 9537
rect 147956 9571 148008 9580
rect 147956 9537 147965 9571
rect 147965 9537 147999 9571
rect 147999 9537 148008 9571
rect 147956 9528 148008 9537
rect 148048 9571 148100 9580
rect 148048 9537 148057 9571
rect 148057 9537 148091 9571
rect 148091 9537 148100 9571
rect 150992 9571 151044 9580
rect 148048 9528 148100 9537
rect 98828 9367 98880 9376
rect 98828 9333 98837 9367
rect 98837 9333 98871 9367
rect 98871 9333 98880 9367
rect 98828 9324 98880 9333
rect 150992 9537 151001 9571
rect 151001 9537 151035 9571
rect 151035 9537 151044 9571
rect 150992 9528 151044 9537
rect 152556 9571 152608 9580
rect 152556 9537 152565 9571
rect 152565 9537 152599 9571
rect 152599 9537 152608 9571
rect 152556 9528 152608 9537
rect 168748 9528 168800 9580
rect 168932 9571 168984 9580
rect 168932 9537 168966 9571
rect 168966 9537 168984 9571
rect 168932 9528 168984 9537
rect 169300 9528 169352 9580
rect 168656 9503 168708 9512
rect 168656 9469 168665 9503
rect 168665 9469 168699 9503
rect 168699 9469 168708 9503
rect 168656 9460 168708 9469
rect 239864 9571 239916 9580
rect 239864 9537 239873 9571
rect 239873 9537 239907 9571
rect 239907 9537 239916 9571
rect 239864 9528 239916 9537
rect 240048 9571 240100 9580
rect 240048 9537 240057 9571
rect 240057 9537 240091 9571
rect 240091 9537 240100 9571
rect 240048 9528 240100 9537
rect 244556 9571 244608 9580
rect 244280 9503 244332 9512
rect 147772 9367 147824 9376
rect 147772 9333 147781 9367
rect 147781 9333 147815 9367
rect 147815 9333 147824 9367
rect 147772 9324 147824 9333
rect 170312 9188 170364 9240
rect 185768 9367 185820 9376
rect 185768 9333 185777 9367
rect 185777 9333 185811 9367
rect 185811 9333 185820 9367
rect 185768 9324 185820 9333
rect 244280 9469 244289 9503
rect 244289 9469 244323 9503
rect 244323 9469 244332 9503
rect 244280 9460 244332 9469
rect 244556 9537 244565 9571
rect 244565 9537 244599 9571
rect 244599 9537 244608 9571
rect 244556 9528 244608 9537
rect 244648 9571 244700 9580
rect 244648 9537 244657 9571
rect 244657 9537 244691 9571
rect 244691 9537 244700 9571
rect 244648 9528 244700 9537
rect 270684 9528 270736 9580
rect 270868 9571 270920 9580
rect 270868 9537 270877 9571
rect 270877 9537 270911 9571
rect 270911 9537 270920 9571
rect 270868 9528 270920 9537
rect 273168 9528 273220 9580
rect 277768 9673 277777 9707
rect 277777 9673 277811 9707
rect 277811 9673 277820 9707
rect 277768 9664 277820 9673
rect 278136 9596 278188 9648
rect 469404 9596 469456 9648
rect 277676 9528 277728 9580
rect 310704 9528 310756 9580
rect 317328 9528 317380 9580
rect 495440 9528 495492 9580
rect 261300 9324 261352 9376
rect 261484 9367 261536 9376
rect 261484 9333 261493 9367
rect 261493 9333 261527 9367
rect 261527 9333 261536 9367
rect 261484 9324 261536 9333
rect 7840 9052 7892 9104
rect 170128 9120 170180 9172
rect 170404 9120 170456 9172
rect 261760 9460 261812 9512
rect 270960 9460 271012 9512
rect 272064 9503 272116 9512
rect 272064 9469 272073 9503
rect 272073 9469 272107 9503
rect 272107 9469 272116 9503
rect 272064 9460 272116 9469
rect 445760 9460 445812 9512
rect 271328 9392 271380 9444
rect 496360 9392 496412 9444
rect 273444 9367 273496 9376
rect 273444 9333 273453 9367
rect 273453 9333 273487 9367
rect 273487 9333 273496 9367
rect 273444 9324 273496 9333
rect 170220 9052 170272 9104
rect 277492 9324 277544 9376
rect 277584 9324 277636 9376
rect 455420 9324 455472 9376
rect 280896 9256 280948 9308
rect 382556 9256 382608 9308
rect 278044 9188 278096 9240
rect 360108 9188 360160 9240
rect 469680 9120 469732 9172
rect 280896 9052 280948 9104
rect 282092 9052 282144 9104
rect 401232 9052 401284 9104
rect 3976 8984 4028 9036
rect 147772 8984 147824 9036
rect 372988 8984 373040 9036
rect 9220 8916 9272 8968
rect 116584 8916 116636 8968
rect 117044 8916 117096 8968
rect 341156 8916 341208 8968
rect 150992 8848 151044 8900
rect 451464 8848 451516 8900
rect 3884 8712 3936 8764
rect 321468 8780 321520 8832
rect 467748 8712 467800 8764
rect 6736 8644 6788 8696
rect 320456 8644 320508 8696
rect 168472 8508 168524 8560
rect 168656 8508 168708 8560
rect 4896 8440 4948 8492
rect 7012 8372 7064 8424
rect 240048 8440 240100 8492
rect 244648 8372 244700 8424
rect 273812 8576 273864 8628
rect 277676 8576 277728 8628
rect 405372 8576 405424 8628
rect 282276 8508 282328 8560
rect 343916 8508 343968 8560
rect 340880 8440 340932 8492
rect 271328 8372 271380 8424
rect 328276 8372 328328 8424
rect 468024 8304 468076 8356
rect 5448 8236 5500 8288
rect 16672 8236 16724 8288
rect 301504 8236 301556 8288
rect 310980 8236 311032 8288
rect 8576 8168 8628 8220
rect 23296 8168 23348 8220
rect 308128 8168 308180 8220
rect 405004 8168 405056 8220
rect 9588 8100 9640 8152
rect 129280 8100 129332 8152
rect 222016 8100 222068 8152
rect 444104 8100 444156 8152
rect 149152 8032 149204 8084
rect 340420 8032 340472 8084
rect 42340 7964 42392 8016
rect 215392 7964 215444 8016
rect 135904 7896 135956 7948
rect 333060 7896 333112 7948
rect 88524 7828 88576 7880
rect 89536 7828 89588 7880
rect 168656 7828 168708 7880
rect 389824 7828 389876 7880
rect 63040 7760 63092 7812
rect 278596 7760 278648 7812
rect 36544 7692 36596 7744
rect 272524 7692 272576 7744
rect 29920 7624 29972 7676
rect 78588 7624 78640 7676
rect 23296 7556 23348 7608
rect 75644 7556 75696 7608
rect 241888 7556 241940 7608
rect 384580 7556 384632 7608
rect 10048 7488 10100 7540
rect 418344 7488 418396 7540
rect 69664 7420 69716 7472
rect 310244 7420 310296 7472
rect 54484 5312 54536 5364
rect 326528 5312 326580 5364
rect 60556 5244 60608 5296
rect 342444 5244 342496 5296
rect 318064 5176 318116 5228
rect 8024 5108 8076 5160
rect 205916 5040 205968 5092
rect 376484 5040 376536 5092
rect 339960 4972 340012 5024
rect 88524 4768 88576 4820
rect 148324 4768 148376 4820
rect 470048 4768 470100 4820
rect 349804 4428 349856 4480
rect 9404 4088 9456 4140
rect 371240 4088 371292 4140
rect 372436 4088 372488 4140
rect 98828 4020 98880 4072
rect 293684 4020 293736 4072
rect 302884 4020 302936 4072
rect 310888 4020 310940 4072
rect 315304 4020 315356 4072
rect 463332 4020 463384 4072
rect 4988 3952 5040 4004
rect 193772 3952 193824 4004
rect 208860 3952 208912 4004
rect 414848 3952 414900 4004
rect 9772 3884 9824 3936
rect 233148 3884 233200 3936
rect 8484 3816 8536 3868
rect 236092 3816 236144 3868
rect 434996 3884 435048 3936
rect 257436 3816 257488 3868
rect 493876 3816 493928 3868
rect 69572 3748 69624 3800
rect 313832 3748 313884 3800
rect 315120 3748 315172 3800
rect 475476 3748 475528 3800
rect 108948 3680 109000 3732
rect 389364 3680 389416 3732
rect 8668 3612 8720 3664
rect 21180 3612 21232 3664
rect 39212 3612 39264 3664
rect 338028 3612 338080 3664
rect 348332 3612 348384 3664
rect 349068 3612 349120 3664
rect 360292 3612 360344 3664
rect 361488 3612 361540 3664
rect 363420 3612 363472 3664
rect 365812 3612 365864 3664
rect 369308 3612 369360 3664
rect 460388 3612 460440 3664
rect 9864 3544 9916 3596
rect 24124 3544 24176 3596
rect 63500 3544 63552 3596
rect 376024 3544 376076 3596
rect 6000 3476 6052 3528
rect 33324 3476 33376 3528
rect 72240 3476 72292 3528
rect 439044 3476 439096 3528
rect 8116 3408 8168 3460
rect 484492 3408 484544 3460
rect 20 3340 72 3392
rect 117044 3340 117096 3392
rect 145380 3340 145432 3392
rect 311256 3340 311308 3392
rect 311900 3340 311952 3392
rect 331864 3340 331916 3392
rect 445116 3340 445168 3392
rect 157340 3272 157392 3324
rect 311992 3272 312044 3324
rect 314384 3272 314436 3324
rect 414940 3272 414992 3324
rect 172612 3204 172664 3256
rect 322296 3204 322348 3256
rect 330484 3204 330536 3256
rect 342260 3204 342312 3256
rect 366364 3204 366416 3256
rect 436100 3204 436152 3256
rect 499764 3204 499816 3256
rect 45284 3136 45336 3188
rect 182180 3136 182232 3188
rect 214932 3136 214984 3188
rect 311348 3136 311400 3188
rect 311440 3136 311492 3188
rect 454316 3136 454368 3188
rect 193772 3068 193824 3120
rect 248420 3068 248472 3120
rect 287612 3068 287664 3120
rect 420552 3068 420604 3120
rect 230204 3000 230256 3052
rect 254308 2932 254360 2984
rect 310520 2932 310572 2984
rect 311164 3000 311216 3052
rect 314844 3000 314896 3052
rect 315948 3000 316000 3052
rect 317972 3000 318024 3052
rect 333520 3000 333572 3052
rect 356796 3000 356848 3052
rect 417884 3000 417936 3052
rect 260380 2864 260432 2916
rect 312636 2864 312688 2916
rect 284668 2796 284720 2848
rect 312084 2796 312136 2848
rect 315580 2932 315632 2984
rect 375564 2932 375616 2984
rect 314292 2864 314344 2916
rect 354220 2864 354272 2916
rect 364248 2864 364300 2916
rect 421012 2864 421064 2916
rect 315764 2796 315816 2848
rect 357348 2796 357400 2848
rect 390652 2796 390704 2848
<< metal2 >>
rect 1646 619520 1758 620960
rect 4590 619520 4702 620960
rect 7718 619520 7830 620960
rect 10662 619520 10774 620960
rect 13606 619520 13718 620960
rect 16734 619520 16846 620960
rect 19678 619520 19790 620960
rect 22806 619520 22918 620960
rect 25750 619520 25862 620960
rect 28878 619520 28990 620960
rect 31822 619520 31934 620960
rect 34950 619520 35062 620960
rect 37894 619520 38006 620960
rect 41022 619520 41134 620960
rect 43966 619520 44078 620960
rect 47094 619520 47206 620960
rect 50038 619520 50150 620960
rect 52982 619520 53094 620960
rect 56110 619520 56222 620960
rect 59054 619520 59166 620960
rect 62182 619520 62294 620960
rect 65126 619520 65238 620960
rect 68254 619520 68366 620960
rect 71198 619520 71310 620960
rect 74326 619520 74438 620960
rect 77270 619520 77382 620960
rect 80398 619520 80510 620960
rect 83342 619520 83454 620960
rect 86470 619520 86582 620960
rect 89414 619520 89526 620960
rect 92358 619520 92470 620960
rect 95486 619520 95598 620960
rect 98430 619520 98542 620960
rect 101558 619520 101670 620960
rect 104502 619520 104614 620960
rect 107630 619520 107742 620960
rect 110574 619520 110686 620960
rect 113702 619520 113814 620960
rect 115952 619534 116532 619562
rect 1688 616146 1716 619520
rect 3422 617808 3478 617817
rect 3422 617743 3478 617752
rect 3436 616894 3464 617743
rect 3424 616888 3476 616894
rect 3424 616830 3476 616836
rect 4632 616758 4660 619520
rect 4620 616752 4672 616758
rect 4620 616694 4672 616700
rect 5448 616752 5500 616758
rect 5448 616694 5500 616700
rect 1676 616140 1728 616146
rect 1676 616082 1728 616088
rect 3054 608832 3110 608841
rect 3054 608767 3056 608776
rect 3108 608767 3110 608776
rect 3056 608738 3108 608744
rect 3424 604512 3476 604518
rect 3422 604480 3424 604489
rect 3476 604480 3478 604489
rect 3422 604415 3478 604424
rect 3514 599856 3570 599865
rect 3514 599791 3570 599800
rect 3528 599350 3556 599791
rect 3516 599344 3568 599350
rect 3516 599286 3568 599292
rect 2778 595504 2834 595513
rect 2778 595439 2834 595448
rect 2792 595066 2820 595439
rect 2780 595060 2832 595066
rect 2780 595002 2832 595008
rect 5172 595060 5224 595066
rect 5172 595002 5224 595008
rect 2780 586560 2832 586566
rect 2778 586528 2780 586537
rect 4896 586560 4948 586566
rect 2832 586528 2834 586537
rect 4896 586502 4948 586508
rect 2778 586463 2834 586472
rect 4804 585608 4856 585614
rect 4804 585550 4856 585556
rect 3608 578400 3660 578406
rect 3608 578342 3660 578348
rect 2778 577552 2834 577561
rect 2778 577487 2834 577496
rect 2792 577318 2820 577487
rect 2780 577312 2832 577318
rect 2780 577254 2832 577260
rect 2870 559600 2926 559609
rect 2870 559535 2926 559544
rect 2884 558958 2912 559535
rect 2872 558952 2924 558958
rect 2872 558894 2924 558900
rect 2778 555248 2834 555257
rect 2778 555183 2834 555192
rect 2792 554810 2820 555183
rect 2780 554804 2832 554810
rect 2780 554746 2832 554752
rect 3146 546272 3202 546281
rect 3146 546207 3202 546216
rect 3160 545154 3188 546207
rect 3148 545148 3200 545154
rect 3148 545090 3200 545096
rect 3424 544264 3476 544270
rect 3424 544206 3476 544212
rect 2870 541648 2926 541657
rect 2870 541583 2926 541592
rect 2884 541006 2912 541583
rect 2872 541000 2924 541006
rect 2872 540942 2924 540948
rect 3146 537296 3202 537305
rect 3146 537231 3202 537240
rect 3160 536858 3188 537231
rect 3148 536852 3200 536858
rect 3148 536794 3200 536800
rect 3330 514992 3386 515001
rect 3330 514927 3386 514936
rect 3344 514826 3372 514927
rect 3332 514820 3384 514826
rect 3332 514762 3384 514768
rect 3146 506016 3202 506025
rect 3146 505951 3202 505960
rect 3160 505170 3188 505951
rect 3148 505164 3200 505170
rect 3148 505106 3200 505112
rect 2778 497040 2834 497049
rect 2778 496975 2780 496984
rect 2832 496975 2834 496984
rect 2780 496946 2832 496952
rect 2778 479088 2834 479097
rect 2778 479023 2780 479032
rect 2832 479023 2834 479032
rect 2780 478994 2832 479000
rect 3330 461136 3386 461145
rect 3330 461071 3386 461080
rect 3344 460970 3372 461071
rect 3332 460964 3384 460970
rect 3332 460906 3384 460912
rect 3146 443184 3202 443193
rect 3146 443119 3202 443128
rect 3056 403232 3108 403238
rect 3056 403174 3108 403180
rect 2962 402928 3018 402937
rect 2962 402863 3018 402872
rect 2976 401674 3004 402863
rect 2964 401668 3016 401674
rect 2964 401610 3016 401616
rect 2778 367024 2834 367033
rect 2778 366959 2834 366968
rect 2792 366722 2820 366959
rect 2780 366716 2832 366722
rect 2780 366658 2832 366664
rect 2964 337544 3016 337550
rect 2964 337486 3016 337492
rect 2872 206032 2924 206038
rect 2870 206000 2872 206009
rect 2924 206000 2926 206009
rect 2870 205935 2926 205944
rect 2780 121168 2832 121174
rect 2780 121110 2832 121116
rect 2792 120873 2820 121110
rect 2778 120864 2834 120873
rect 2778 120799 2834 120808
rect 2976 101114 3004 337486
rect 3068 317801 3096 403174
rect 3160 336734 3188 443119
rect 3330 434208 3386 434217
rect 3330 434143 3386 434152
rect 3344 433362 3372 434143
rect 3332 433356 3384 433362
rect 3332 433298 3384 433304
rect 3238 429856 3294 429865
rect 3238 429791 3294 429800
rect 3148 336728 3200 336734
rect 3148 336670 3200 336676
rect 3054 317792 3110 317801
rect 3054 317727 3110 317736
rect 3252 273358 3280 429791
rect 3330 425232 3386 425241
rect 3330 425167 3332 425176
rect 3384 425167 3386 425176
rect 3332 425138 3384 425144
rect 3330 407280 3386 407289
rect 3330 407215 3386 407224
rect 3344 407182 3372 407215
rect 3332 407176 3384 407182
rect 3332 407118 3384 407124
rect 3332 407040 3384 407046
rect 3332 406982 3384 406988
rect 3240 273352 3292 273358
rect 3240 273294 3292 273300
rect 3240 252748 3292 252754
rect 3240 252690 3292 252696
rect 3054 223952 3110 223961
rect 3054 223887 3110 223896
rect 3068 223786 3096 223887
rect 3056 223780 3108 223786
rect 3056 223722 3108 223728
rect 3252 201385 3280 252690
rect 3344 246265 3372 406982
rect 3330 246256 3386 246265
rect 3330 246191 3386 246200
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 3238 201376 3294 201385
rect 3238 201311 3294 201320
rect 3240 197804 3292 197810
rect 3240 197746 3292 197752
rect 3056 183456 3108 183462
rect 3054 183424 3056 183433
rect 3108 183424 3110 183433
rect 3054 183359 3110 183368
rect 3148 157072 3200 157078
rect 3148 157014 3200 157020
rect 3160 156777 3188 157014
rect 3146 156768 3202 156777
rect 3146 156703 3202 156712
rect 3146 117328 3202 117337
rect 3146 117263 3202 117272
rect 2964 101108 3016 101114
rect 2964 101050 3016 101056
rect 2780 76968 2832 76974
rect 2780 76910 2832 76916
rect 2792 75993 2820 76910
rect 2778 75984 2834 75993
rect 2778 75919 2834 75928
rect 3160 67017 3188 117263
rect 3146 67008 3202 67017
rect 3146 66943 3202 66952
rect 2780 58268 2832 58274
rect 2780 58210 2832 58216
rect 2792 58041 2820 58210
rect 2778 58032 2834 58041
rect 2778 57967 2834 57976
rect 2780 53712 2832 53718
rect 2778 53680 2780 53689
rect 2832 53680 2834 53689
rect 2778 53615 2834 53624
rect 3252 40361 3280 197746
rect 3344 188057 3372 222527
rect 3330 188048 3386 188057
rect 3330 187983 3386 187992
rect 3330 179072 3386 179081
rect 3330 179007 3386 179016
rect 3344 178906 3372 179007
rect 3332 178900 3384 178906
rect 3332 178842 3384 178848
rect 3344 170202 3372 178842
rect 3332 170196 3384 170202
rect 3332 170138 3384 170144
rect 3332 161152 3384 161158
rect 3330 161120 3332 161129
rect 3384 161120 3386 161129
rect 3330 161055 3386 161064
rect 3332 138984 3384 138990
rect 3332 138926 3384 138932
rect 3344 138825 3372 138926
rect 3330 138816 3386 138825
rect 3330 138751 3386 138760
rect 3332 100768 3384 100774
rect 3332 100710 3384 100716
rect 3238 40352 3294 40361
rect 3238 40287 3294 40296
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8809 2820 9318
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 3344 8673 3372 100710
rect 3436 35737 3464 544206
rect 3516 536648 3568 536654
rect 3516 536590 3568 536596
rect 3528 80617 3556 536590
rect 3620 389706 3648 578342
rect 4528 533792 4580 533798
rect 4528 533734 4580 533740
rect 3698 528320 3754 528329
rect 3698 528255 3754 528264
rect 3712 494222 3740 528255
rect 3882 519344 3938 519353
rect 3882 519279 3938 519288
rect 3700 494216 3752 494222
rect 3700 494158 3752 494164
rect 3698 420880 3754 420889
rect 3698 420815 3754 420824
rect 3608 389700 3660 389706
rect 3608 389642 3660 389648
rect 3606 389600 3662 389609
rect 3606 389535 3662 389544
rect 3620 389230 3648 389535
rect 3608 389224 3660 389230
rect 3608 389166 3660 389172
rect 3608 332580 3660 332586
rect 3608 332522 3660 332528
rect 3620 331401 3648 332522
rect 3606 331392 3662 331401
rect 3606 331327 3662 331336
rect 3606 322416 3662 322425
rect 3606 322351 3662 322360
rect 3620 321638 3648 322351
rect 3608 321632 3660 321638
rect 3608 321574 3660 321580
rect 3606 290864 3662 290873
rect 3606 290799 3662 290808
rect 3620 289882 3648 290799
rect 3608 289876 3660 289882
rect 3608 289818 3660 289824
rect 3608 273216 3660 273222
rect 3606 273184 3608 273193
rect 3660 273184 3662 273193
rect 3606 273119 3662 273128
rect 3606 268560 3662 268569
rect 3606 268495 3662 268504
rect 3620 267782 3648 268495
rect 3608 267776 3660 267782
rect 3608 267718 3660 267724
rect 3608 219428 3660 219434
rect 3608 219370 3660 219376
rect 3620 219337 3648 219370
rect 3606 219328 3662 219337
rect 3606 219263 3662 219272
rect 3608 217660 3660 217666
rect 3608 217602 3660 217608
rect 3620 214985 3648 217602
rect 3606 214976 3662 214985
rect 3606 214911 3662 214920
rect 3712 118454 3740 420815
rect 3790 416256 3846 416265
rect 3790 416191 3846 416200
rect 3804 395622 3832 416191
rect 3792 395616 3844 395622
rect 3792 395558 3844 395564
rect 3792 389700 3844 389706
rect 3792 389642 3844 389648
rect 3804 384985 3832 389642
rect 3790 384976 3846 384985
rect 3790 384911 3846 384920
rect 3792 356108 3844 356114
rect 3792 356050 3844 356056
rect 3700 118448 3752 118454
rect 3700 118390 3752 118396
rect 3698 118008 3754 118017
rect 3698 117943 3754 117952
rect 3712 101114 3740 117943
rect 3700 101108 3752 101114
rect 3700 101050 3752 101056
rect 3804 84969 3832 356050
rect 3896 304774 3924 519279
rect 3976 417580 4028 417586
rect 3976 417522 4028 417528
rect 3884 304768 3936 304774
rect 3884 304710 3936 304716
rect 3884 298376 3936 298382
rect 3884 298318 3936 298324
rect 3896 264217 3924 298318
rect 3882 264208 3938 264217
rect 3882 264143 3938 264152
rect 3882 255232 3938 255241
rect 3882 255167 3938 255176
rect 3790 84960 3846 84969
rect 3790 84895 3846 84904
rect 3514 80608 3570 80617
rect 3514 80543 3570 80552
rect 3422 35728 3478 35737
rect 3422 35663 3478 35672
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 3330 8664 3386 8673
rect 3330 8599 3386 8608
rect 3436 7993 3464 17711
rect 3896 8770 3924 255167
rect 3988 178906 4016 417522
rect 4068 411528 4120 411534
rect 4068 411470 4120 411476
rect 4080 407046 4108 411470
rect 4068 407040 4120 407046
rect 4068 406982 4120 406988
rect 4068 335776 4120 335782
rect 4068 335718 4120 335724
rect 3976 178900 4028 178906
rect 3976 178842 4028 178848
rect 3976 169856 4028 169862
rect 3976 169798 4028 169804
rect 3988 143177 4016 169798
rect 4080 152153 4108 335718
rect 4158 308816 4214 308825
rect 4158 308751 4214 308760
rect 4172 303142 4200 308751
rect 4160 303136 4212 303142
rect 4160 303078 4212 303084
rect 4436 219496 4488 219502
rect 4436 219438 4488 219444
rect 4066 152144 4122 152153
rect 4066 152079 4122 152088
rect 3974 143168 4030 143177
rect 3974 143103 4030 143112
rect 3988 125594 4016 143103
rect 4448 142154 4476 219438
rect 4172 142126 4476 142154
rect 4066 134192 4122 134201
rect 4172 134178 4200 142126
rect 4122 134150 4200 134178
rect 4066 134127 4122 134136
rect 4066 129840 4122 129849
rect 4066 129775 4122 129784
rect 3976 125588 4028 125594
rect 3976 125530 4028 125536
rect 3974 125216 4030 125225
rect 3974 125151 4030 125160
rect 3988 9042 4016 125151
rect 4080 121854 4108 129775
rect 4540 127566 4568 533734
rect 4712 366716 4764 366722
rect 4712 366658 4764 366664
rect 4620 348288 4672 348294
rect 4620 348230 4672 348236
rect 4632 251122 4660 348230
rect 4724 325582 4752 366658
rect 4712 325576 4764 325582
rect 4712 325518 4764 325524
rect 4712 304224 4764 304230
rect 4712 304166 4764 304172
rect 4620 251116 4672 251122
rect 4620 251058 4672 251064
rect 4620 218952 4672 218958
rect 4620 218894 4672 218900
rect 4528 127560 4580 127566
rect 4528 127502 4580 127508
rect 4068 121848 4120 121854
rect 4068 121790 4120 121796
rect 4632 118590 4660 218894
rect 4620 118584 4672 118590
rect 4620 118526 4672 118532
rect 4066 111888 4122 111897
rect 4066 111823 4122 111832
rect 4080 44713 4108 111823
rect 4724 76974 4752 304166
rect 4712 76968 4764 76974
rect 4712 76910 4764 76916
rect 4066 44704 4122 44713
rect 4066 44639 4122 44648
rect 4816 9382 4844 585550
rect 4908 118998 4936 586502
rect 4988 577312 5040 577318
rect 4988 577254 5040 577260
rect 4896 118992 4948 118998
rect 4896 118934 4948 118940
rect 4896 118448 4948 118454
rect 4896 118390 4948 118396
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8764 3936 8770
rect 3884 8706 3936 8712
rect 4908 8498 4936 118390
rect 5000 110566 5028 577254
rect 5080 417376 5132 417382
rect 5080 417318 5132 417324
rect 5092 169998 5120 417318
rect 5184 327758 5212 595002
rect 5356 497004 5408 497010
rect 5356 496946 5408 496952
rect 5264 479052 5316 479058
rect 5264 478994 5316 479000
rect 5276 344486 5304 478994
rect 5368 375630 5396 496946
rect 5356 375624 5408 375630
rect 5356 375566 5408 375572
rect 5264 344480 5316 344486
rect 5264 344422 5316 344428
rect 5356 336728 5408 336734
rect 5356 336670 5408 336676
rect 5264 329044 5316 329050
rect 5264 328986 5316 328992
rect 5172 327752 5224 327758
rect 5172 327694 5224 327700
rect 5172 236360 5224 236366
rect 5172 236302 5224 236308
rect 5184 170066 5212 236302
rect 5172 170060 5224 170066
rect 5172 170002 5224 170008
rect 5080 169992 5132 169998
rect 5080 169934 5132 169940
rect 5080 127424 5132 127430
rect 5080 127366 5132 127372
rect 5092 113174 5120 127366
rect 5276 121174 5304 328986
rect 5368 129878 5396 336670
rect 5460 220153 5488 616694
rect 6828 616276 6880 616282
rect 6828 616218 6880 616224
rect 6184 608796 6236 608802
rect 6184 608738 6236 608744
rect 5908 475584 5960 475590
rect 5908 475526 5960 475532
rect 5816 304768 5868 304774
rect 5816 304710 5868 304716
rect 5632 281376 5684 281382
rect 5632 281318 5684 281324
rect 5446 220144 5502 220153
rect 5446 220079 5502 220088
rect 5448 219020 5500 219026
rect 5448 218962 5500 218968
rect 5356 129872 5408 129878
rect 5356 129814 5408 129820
rect 5356 125588 5408 125594
rect 5356 125530 5408 125536
rect 5264 121168 5316 121174
rect 5264 121110 5316 121116
rect 5092 113146 5304 113174
rect 5276 110838 5304 113146
rect 5264 110832 5316 110838
rect 5264 110774 5316 110780
rect 4988 110560 5040 110566
rect 4988 110502 5040 110508
rect 5080 108588 5132 108594
rect 5080 108530 5132 108536
rect 4988 100836 5040 100842
rect 4988 100778 5040 100784
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 3422 7984 3478 7993
rect 3422 7919 3478 7928
rect 5000 4010 5028 100778
rect 5092 53718 5120 108530
rect 5172 108316 5224 108322
rect 5172 108258 5224 108264
rect 5184 58274 5212 108258
rect 5276 100774 5304 110774
rect 5264 100768 5316 100774
rect 5264 100710 5316 100716
rect 5368 89690 5396 125530
rect 5356 89684 5408 89690
rect 5356 89626 5408 89632
rect 5172 58268 5224 58274
rect 5172 58210 5224 58216
rect 5080 53712 5132 53718
rect 5080 53654 5132 53660
rect 5460 8294 5488 218962
rect 5644 206038 5672 281318
rect 5724 218544 5776 218550
rect 5724 218486 5776 218492
rect 5632 206032 5684 206038
rect 5632 205974 5684 205980
rect 5632 203720 5684 203726
rect 5632 203662 5684 203668
rect 5644 111382 5672 203662
rect 5736 120018 5764 218486
rect 5724 120012 5776 120018
rect 5724 119954 5776 119960
rect 5828 118289 5856 304710
rect 5920 304570 5948 475526
rect 6092 393440 6144 393446
rect 6092 393382 6144 393388
rect 5908 304564 5960 304570
rect 5908 304506 5960 304512
rect 5908 223780 5960 223786
rect 5908 223722 5960 223728
rect 5920 119270 5948 223722
rect 6000 209568 6052 209574
rect 6000 209510 6052 209516
rect 5908 119264 5960 119270
rect 5908 119206 5960 119212
rect 5814 118280 5870 118289
rect 5814 118215 5870 118224
rect 5632 111376 5684 111382
rect 5632 111318 5684 111324
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 6012 3534 6040 209510
rect 6104 183462 6132 393382
rect 6092 183456 6144 183462
rect 6092 183398 6144 183404
rect 6196 117706 6224 608738
rect 6276 554804 6328 554810
rect 6276 554746 6328 554752
rect 6288 118318 6316 554746
rect 6368 537736 6420 537742
rect 6368 537678 6420 537684
rect 6380 157078 6408 537678
rect 6736 536852 6788 536858
rect 6736 536794 6788 536800
rect 6460 494624 6512 494630
rect 6460 494566 6512 494572
rect 6472 161158 6500 494566
rect 6552 463072 6604 463078
rect 6552 463014 6604 463020
rect 6460 161152 6512 161158
rect 6460 161094 6512 161100
rect 6368 157072 6420 157078
rect 6368 157014 6420 157020
rect 6564 138990 6592 463014
rect 6644 425196 6696 425202
rect 6644 425138 6696 425144
rect 6552 138984 6604 138990
rect 6552 138926 6604 138932
rect 6276 118312 6328 118318
rect 6276 118254 6328 118260
rect 6184 117700 6236 117706
rect 6184 117642 6236 117648
rect 6656 111246 6684 425138
rect 6748 265742 6776 536794
rect 6736 265736 6788 265742
rect 6736 265678 6788 265684
rect 6736 218612 6788 218618
rect 6736 218554 6788 218560
rect 6644 111240 6696 111246
rect 6644 111182 6696 111188
rect 6184 100768 6236 100774
rect 6184 100710 6236 100716
rect 6196 79762 6224 100710
rect 6184 79756 6236 79762
rect 6184 79698 6236 79704
rect 6748 8702 6776 218554
rect 6840 110634 6868 616218
rect 9864 616208 9916 616214
rect 9864 616150 9916 616156
rect 7840 513732 7892 513738
rect 7840 513674 7892 513680
rect 7104 487212 7156 487218
rect 7104 487154 7156 487160
rect 6920 218680 6972 218686
rect 6920 218622 6972 218628
rect 6932 149161 6960 218622
rect 7010 158808 7066 158817
rect 7010 158743 7066 158752
rect 6918 149152 6974 149161
rect 6918 149087 6974 149096
rect 7024 120154 7052 158743
rect 7116 120630 7144 487154
rect 7564 311908 7616 311914
rect 7564 311850 7616 311856
rect 7196 222284 7248 222290
rect 7196 222226 7248 222232
rect 7208 120834 7236 222226
rect 7288 218476 7340 218482
rect 7288 218418 7340 218424
rect 7196 120828 7248 120834
rect 7196 120770 7248 120776
rect 7104 120624 7156 120630
rect 7104 120566 7156 120572
rect 7012 120148 7064 120154
rect 7012 120090 7064 120096
rect 7024 113174 7052 120090
rect 7300 113937 7328 218418
rect 7472 217524 7524 217530
rect 7472 217466 7524 217472
rect 7378 197840 7434 197849
rect 7378 197775 7434 197784
rect 7392 169862 7420 197775
rect 7484 178945 7512 217466
rect 7576 197810 7604 311850
rect 7852 300150 7880 513674
rect 8024 509312 8076 509318
rect 8024 509254 8076 509260
rect 7932 343936 7984 343942
rect 7932 343878 7984 343884
rect 7840 300144 7892 300150
rect 7840 300086 7892 300092
rect 7852 296714 7880 300086
rect 7668 296686 7880 296714
rect 7564 197804 7616 197810
rect 7564 197746 7616 197752
rect 7470 178936 7526 178945
rect 7470 178871 7526 178880
rect 7380 169856 7432 169862
rect 7380 169798 7432 169804
rect 7378 168464 7434 168473
rect 7378 168399 7434 168408
rect 7286 113928 7342 113937
rect 7286 113863 7342 113872
rect 7024 113146 7236 113174
rect 6828 110628 6880 110634
rect 6828 110570 6880 110576
rect 7012 109200 7064 109206
rect 7012 109142 7064 109148
rect 6736 8696 6788 8702
rect 6736 8638 6788 8644
rect 7024 8430 7052 109142
rect 7104 108384 7156 108390
rect 7104 108326 7156 108332
rect 7116 58546 7144 108326
rect 7104 58540 7156 58546
rect 7104 58482 7156 58488
rect 7208 49609 7236 113146
rect 7392 59265 7420 168399
rect 7484 68921 7512 178871
rect 7562 149152 7618 149161
rect 7562 149087 7618 149096
rect 7470 68912 7526 68921
rect 7470 68847 7526 68856
rect 7378 59256 7434 59265
rect 7378 59191 7434 59200
rect 7194 49600 7250 49609
rect 7194 49535 7250 49544
rect 7576 39953 7604 149087
rect 7668 139777 7696 296686
rect 7840 219360 7892 219366
rect 7840 219302 7892 219308
rect 7748 219292 7800 219298
rect 7748 219234 7800 219240
rect 7654 139768 7710 139777
rect 7654 139703 7710 139712
rect 7562 39944 7618 39953
rect 7562 39879 7618 39888
rect 7668 30297 7696 139703
rect 7654 30288 7710 30297
rect 7654 30223 7710 30232
rect 7760 9450 7788 219234
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7852 9110 7880 219302
rect 7944 108633 7972 343878
rect 8036 208321 8064 509254
rect 9588 487280 9640 487286
rect 9588 487222 9640 487228
rect 8944 469600 8996 469606
rect 8944 469542 8996 469548
rect 8116 415336 8168 415342
rect 8116 415278 8168 415284
rect 8022 208312 8078 208321
rect 8022 208247 8078 208256
rect 7930 108624 7986 108633
rect 7930 108559 7986 108568
rect 8036 98841 8064 208247
rect 8022 98832 8078 98841
rect 8022 98767 8078 98776
rect 8024 89684 8076 89690
rect 8024 89626 8076 89632
rect 8036 89049 8064 89626
rect 8022 89040 8078 89049
rect 8022 88975 8078 88984
rect 8128 78577 8156 415278
rect 8852 375556 8904 375562
rect 8852 375498 8904 375504
rect 8300 295656 8352 295662
rect 8300 295598 8352 295604
rect 8208 219156 8260 219162
rect 8208 219098 8260 219104
rect 8220 189009 8248 219098
rect 8206 189000 8262 189009
rect 8206 188935 8262 188944
rect 8206 129976 8262 129985
rect 8206 129911 8262 129920
rect 8220 129878 8248 129911
rect 8208 129872 8260 129878
rect 8208 129814 8260 129820
rect 8114 78568 8170 78577
rect 8114 78503 8170 78512
rect 8114 59256 8170 59265
rect 8114 59191 8170 59200
rect 8024 42152 8076 42158
rect 8024 42094 8076 42100
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 8036 5166 8064 42094
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 8128 3466 8156 59191
rect 8220 20505 8248 129814
rect 8312 79626 8340 295598
rect 8484 219224 8536 219230
rect 8484 219166 8536 219172
rect 8392 217592 8444 217598
rect 8392 217534 8444 217540
rect 8404 136474 8432 217534
rect 8392 136468 8444 136474
rect 8392 136410 8444 136416
rect 8496 136270 8524 219166
rect 8576 218884 8628 218890
rect 8576 218826 8628 218832
rect 8484 136264 8536 136270
rect 8484 136206 8536 136212
rect 8588 133142 8616 218826
rect 8760 218816 8812 218822
rect 8760 218758 8812 218764
rect 8668 203924 8720 203930
rect 8668 203866 8720 203872
rect 8576 133136 8628 133142
rect 8576 133078 8628 133084
rect 8576 109744 8628 109750
rect 8576 109686 8628 109692
rect 8484 109336 8536 109342
rect 8484 109278 8536 109284
rect 8392 108452 8444 108458
rect 8392 108394 8444 108400
rect 8300 79620 8352 79626
rect 8300 79562 8352 79568
rect 8404 42294 8432 108394
rect 8392 42288 8444 42294
rect 8392 42230 8444 42236
rect 8206 20496 8262 20505
rect 8206 20431 8262 20440
rect 8496 3874 8524 109278
rect 8588 8226 8616 109686
rect 8680 109206 8708 203866
rect 8668 109200 8720 109206
rect 8668 109142 8720 109148
rect 8668 109064 8720 109070
rect 8668 109006 8720 109012
rect 8576 8220 8628 8226
rect 8576 8162 8628 8168
rect 8484 3868 8536 3874
rect 8484 3810 8536 3816
rect 8680 3670 8708 109006
rect 8772 9586 8800 218758
rect 8864 79898 8892 375498
rect 8956 156942 8984 469542
rect 9404 349376 9456 349382
rect 9404 349318 9456 349324
rect 9128 333056 9180 333062
rect 9128 332998 9180 333004
rect 9140 332858 9168 332998
rect 9128 332852 9180 332858
rect 9128 332794 9180 332800
rect 9036 263968 9088 263974
rect 9036 263910 9088 263916
rect 8944 156936 8996 156942
rect 8944 156878 8996 156884
rect 8944 136264 8996 136270
rect 8944 136206 8996 136212
rect 8956 121417 8984 136206
rect 9048 133074 9076 263910
rect 9140 157146 9168 332794
rect 9220 324896 9272 324902
rect 9220 324838 9272 324844
rect 9128 157140 9180 157146
rect 9128 157082 9180 157088
rect 9128 136468 9180 136474
rect 9128 136410 9180 136416
rect 9036 133068 9088 133074
rect 9036 133010 9088 133016
rect 9140 132954 9168 136410
rect 9232 133074 9260 324838
rect 9312 252680 9364 252686
rect 9312 252622 9364 252628
rect 9220 133068 9272 133074
rect 9220 133010 9272 133016
rect 9140 132926 9260 132954
rect 9128 132864 9180 132870
rect 9128 132806 9180 132812
rect 9140 121922 9168 132806
rect 9128 121916 9180 121922
rect 9128 121858 9180 121864
rect 8942 121408 8998 121417
rect 8942 121343 8998 121352
rect 9036 111580 9088 111586
rect 9036 111522 9088 111528
rect 8944 108520 8996 108526
rect 8944 108462 8996 108468
rect 8852 79892 8904 79898
rect 8852 79834 8904 79840
rect 8956 79694 8984 108462
rect 8944 79688 8996 79694
rect 8944 79630 8996 79636
rect 9048 66026 9076 111522
rect 9126 109168 9182 109177
rect 9126 109103 9182 109112
rect 9140 79830 9168 109103
rect 9128 79824 9180 79830
rect 9128 79766 9180 79772
rect 9128 79688 9180 79694
rect 9128 79630 9180 79636
rect 9036 66020 9088 66026
rect 9036 65962 9088 65968
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 9140 9489 9168 79630
rect 9232 66162 9260 132926
rect 9220 66156 9272 66162
rect 9220 66098 9272 66104
rect 9324 25906 9352 252622
rect 9416 133074 9444 349318
rect 9496 218748 9548 218754
rect 9496 218690 9548 218696
rect 9508 217841 9536 218690
rect 9494 217832 9550 217841
rect 9494 217767 9550 217776
rect 9496 217728 9548 217734
rect 9496 217670 9548 217676
rect 9508 203930 9536 217670
rect 9496 203924 9548 203930
rect 9496 203866 9548 203872
rect 9404 133068 9456 133074
rect 9404 133010 9456 133016
rect 9496 133000 9548 133006
rect 9496 132942 9548 132948
rect 9404 132932 9456 132938
rect 9404 132874 9456 132880
rect 9416 54874 9444 132874
rect 9508 121786 9536 132942
rect 9496 121780 9548 121786
rect 9496 121722 9548 121728
rect 9496 107704 9548 107710
rect 9496 107646 9548 107652
rect 9508 101046 9536 107646
rect 9496 101040 9548 101046
rect 9496 100982 9548 100988
rect 9404 54868 9456 54874
rect 9404 54810 9456 54816
rect 9404 42016 9456 42022
rect 9404 41958 9456 41964
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9232 8974 9260 25638
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9416 4146 9444 41958
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9508 11898 9536 25774
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9600 8158 9628 487222
rect 9772 475380 9824 475386
rect 9772 475322 9824 475328
rect 9680 422612 9732 422618
rect 9680 422554 9732 422560
rect 9692 118658 9720 422554
rect 9784 142322 9812 475322
rect 9772 142316 9824 142322
rect 9772 142258 9824 142264
rect 9772 142180 9824 142186
rect 9772 142122 9824 142128
rect 9680 118652 9732 118658
rect 9680 118594 9732 118600
rect 9588 8152 9640 8158
rect 9588 8094 9640 8100
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9784 3942 9812 142122
rect 9876 132938 9904 616150
rect 13648 615494 13676 619520
rect 22848 616826 22876 619520
rect 22836 616820 22888 616826
rect 22836 616762 22888 616768
rect 23388 616820 23440 616826
rect 23388 616762 23440 616768
rect 17224 616480 17276 616486
rect 17224 616422 17276 616428
rect 13648 615466 13768 615494
rect 12992 527944 13044 527950
rect 12992 527886 13044 527892
rect 12716 527876 12768 527882
rect 12716 527818 12768 527824
rect 11428 524544 11480 524550
rect 11428 524486 11480 524492
rect 11440 304842 11468 524486
rect 12728 518894 12756 527818
rect 12728 518866 12848 518894
rect 11704 407176 11756 407182
rect 11704 407118 11756 407124
rect 11716 317286 11744 407118
rect 11796 395208 11848 395214
rect 11796 395150 11848 395156
rect 11704 317280 11756 317286
rect 11704 317222 11756 317228
rect 11428 304836 11480 304842
rect 11428 304778 11480 304784
rect 11808 219570 11836 395150
rect 12820 219570 12848 518866
rect 13004 249830 13032 527886
rect 13740 383246 13768 615466
rect 15016 561740 15068 561746
rect 15016 561682 15068 561688
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 13728 383240 13780 383246
rect 13728 383182 13780 383188
rect 14476 326670 14504 514762
rect 15028 423570 15056 561682
rect 15292 561672 15344 561678
rect 15292 561614 15344 561620
rect 15304 525094 15332 561614
rect 15292 525088 15344 525094
rect 15292 525030 15344 525036
rect 16212 480480 16264 480486
rect 16212 480422 16264 480428
rect 15016 423564 15068 423570
rect 15016 423506 15068 423512
rect 14464 326664 14516 326670
rect 14464 326606 14516 326612
rect 12992 249824 13044 249830
rect 12992 249766 13044 249772
rect 15568 222216 15620 222222
rect 15568 222158 15620 222164
rect 15580 219994 15608 222158
rect 15226 219966 15608 219994
rect 16224 219570 16252 480422
rect 17236 219570 17264 616422
rect 23020 600772 23072 600778
rect 23020 600714 23072 600720
rect 21640 487348 21692 487354
rect 21640 487290 21692 487296
rect 21652 306066 21680 487290
rect 22836 480684 22888 480690
rect 22836 480626 22888 480632
rect 22848 394874 22876 480626
rect 22836 394868 22888 394874
rect 22836 394810 22888 394816
rect 22928 394732 22980 394738
rect 22928 394674 22980 394680
rect 22100 387048 22152 387054
rect 22100 386990 22152 386996
rect 22112 306202 22140 386990
rect 22100 306196 22152 306202
rect 22100 306138 22152 306144
rect 21640 306060 21692 306066
rect 21640 306002 21692 306008
rect 21548 305856 21600 305862
rect 21548 305798 21600 305804
rect 20536 237584 20588 237590
rect 20536 237526 20588 237532
rect 11796 219564 11848 219570
rect 11796 219506 11848 219512
rect 12808 219564 12860 219570
rect 12808 219506 12860 219512
rect 16212 219564 16264 219570
rect 16212 219506 16264 219512
rect 17224 219564 17276 219570
rect 17224 219506 17276 219512
rect 20548 219366 20576 237526
rect 21560 219366 21588 305798
rect 21640 222284 21692 222290
rect 21640 222226 21692 222232
rect 21652 219994 21680 222226
rect 21652 219966 21850 219994
rect 22940 219366 22968 394674
rect 23032 220114 23060 600714
rect 23400 310758 23428 616762
rect 25792 616214 25820 619520
rect 28920 616214 28948 619520
rect 34992 616826 35020 619520
rect 34980 616820 35032 616826
rect 34980 616762 35032 616768
rect 35808 616820 35860 616826
rect 35808 616762 35860 616768
rect 25780 616208 25832 616214
rect 25780 616150 25832 616156
rect 28908 616208 28960 616214
rect 28908 616150 28960 616156
rect 28908 580780 28960 580786
rect 28908 580722 28960 580728
rect 27436 524612 27488 524618
rect 27436 524554 27488 524560
rect 27448 423026 27476 524554
rect 27528 489524 27580 489530
rect 27528 489466 27580 489472
rect 27540 423162 27568 489466
rect 27528 423156 27580 423162
rect 27528 423098 27580 423104
rect 27436 423020 27488 423026
rect 27436 422962 27488 422968
rect 23388 310752 23440 310758
rect 23388 310694 23440 310700
rect 23020 220108 23072 220114
rect 23020 220050 23072 220056
rect 28920 219994 28948 580722
rect 29644 493196 29696 493202
rect 29644 493138 29696 493144
rect 29656 487082 29684 493138
rect 32310 493096 32366 493105
rect 32310 493031 32312 493040
rect 32364 493031 32366 493040
rect 32312 493002 32364 493008
rect 32404 492992 32456 492998
rect 32404 492934 32456 492940
rect 32772 492992 32824 492998
rect 32772 492934 32824 492940
rect 32416 492697 32444 492934
rect 32402 492688 32458 492697
rect 32402 492623 32458 492632
rect 29644 487076 29696 487082
rect 29644 487018 29696 487024
rect 32784 224262 32812 492934
rect 35820 406094 35848 616762
rect 36360 616548 36412 616554
rect 36360 616490 36412 616496
rect 35808 406088 35860 406094
rect 35808 406030 35860 406036
rect 36372 266354 36400 616490
rect 44008 615494 44036 619520
rect 53024 616826 53052 619520
rect 53012 616820 53064 616826
rect 53012 616762 53064 616768
rect 53748 616820 53800 616826
rect 53748 616762 53800 616768
rect 44008 615466 44128 615494
rect 43076 572756 43128 572762
rect 43076 572698 43128 572704
rect 41788 507204 41840 507210
rect 41788 507146 41840 507152
rect 41800 439346 41828 507146
rect 41788 439340 41840 439346
rect 41788 439282 41840 439288
rect 43088 395826 43116 572698
rect 43168 451308 43220 451314
rect 43168 451250 43220 451256
rect 43180 439482 43208 451250
rect 43168 439476 43220 439482
rect 43168 439418 43220 439424
rect 44100 434926 44128 615466
rect 50160 599072 50212 599078
rect 50158 599040 50160 599049
rect 50212 599040 50214 599049
rect 50158 598975 50214 598984
rect 51448 561740 51500 561746
rect 51448 561682 51500 561688
rect 46020 513800 46072 513806
rect 46020 513742 46072 513748
rect 45744 513664 45796 513670
rect 45744 513606 45796 513612
rect 44088 434920 44140 434926
rect 44088 434862 44140 434868
rect 43076 395820 43128 395826
rect 43076 395762 43128 395768
rect 45756 394806 45784 513606
rect 46032 424522 46060 513742
rect 46204 513732 46256 513738
rect 46204 513674 46256 513680
rect 46020 424516 46072 424522
rect 46020 424458 46072 424464
rect 45744 394800 45796 394806
rect 45744 394742 45796 394748
rect 39408 381070 39436 381101
rect 39396 381064 39448 381070
rect 39394 381032 39396 381041
rect 39448 381032 39450 381041
rect 39394 380967 39450 380976
rect 39408 380934 39436 380967
rect 39396 380928 39448 380934
rect 39396 380870 39448 380876
rect 40592 380928 40644 380934
rect 40592 380870 40644 380876
rect 38842 333296 38898 333305
rect 38842 333231 38844 333240
rect 38896 333231 38898 333240
rect 38844 333202 38896 333208
rect 36360 266348 36412 266354
rect 36360 266290 36412 266296
rect 40604 226982 40632 380870
rect 46216 329254 46244 513674
rect 47676 435056 47728 435062
rect 47674 435024 47676 435033
rect 47728 435024 47730 435033
rect 47674 434959 47730 434968
rect 48044 434988 48096 434994
rect 48044 434930 48096 434936
rect 48228 434988 48280 434994
rect 48228 434930 48280 434936
rect 47860 434852 47912 434858
rect 47860 434794 47912 434800
rect 47872 434602 47900 434794
rect 48056 434761 48084 434930
rect 48136 434920 48188 434926
rect 48136 434862 48188 434868
rect 48042 434752 48098 434761
rect 48042 434687 48098 434696
rect 48148 434602 48176 434862
rect 47872 434574 48176 434602
rect 48240 329322 48268 434930
rect 48228 329316 48280 329322
rect 48228 329258 48280 329264
rect 46204 329248 46256 329254
rect 46204 329190 46256 329196
rect 51460 304774 51488 561682
rect 53472 451104 53524 451110
rect 53472 451046 53524 451052
rect 53484 446962 53512 451046
rect 53472 446956 53524 446962
rect 53472 446898 53524 446904
rect 51448 304768 51500 304774
rect 51448 304710 51500 304716
rect 40592 226976 40644 226982
rect 40592 226918 40644 226924
rect 32772 224256 32824 224262
rect 32772 224198 32824 224204
rect 42064 223372 42116 223378
rect 42064 223314 42116 223320
rect 35164 222964 35216 222970
rect 35164 222906 35216 222912
rect 28474 219966 28948 219994
rect 34794 220008 34850 220017
rect 35176 219994 35204 222906
rect 42076 220017 42104 223314
rect 48688 222284 48740 222290
rect 48688 222226 48740 222232
rect 42062 220008 42118 220017
rect 34850 219966 35204 219994
rect 41722 219966 42062 219994
rect 34794 219943 34850 219952
rect 48700 219994 48728 222226
rect 49976 220448 50028 220454
rect 49976 220390 50028 220396
rect 49988 220017 50016 220390
rect 48346 219966 48728 219994
rect 49974 220008 50030 220017
rect 42062 219943 42118 219952
rect 49974 219943 50030 219952
rect 42076 219883 42104 219943
rect 53760 219502 53788 616762
rect 65168 616758 65196 619520
rect 65156 616752 65208 616758
rect 65156 616694 65208 616700
rect 66168 616752 66220 616758
rect 66168 616694 66220 616700
rect 55496 604512 55548 604518
rect 55496 604454 55548 604460
rect 53840 599412 53892 599418
rect 53840 599354 53892 599360
rect 53852 222698 53880 599354
rect 54024 451308 54076 451314
rect 54024 451250 54076 451256
rect 53932 451104 53984 451110
rect 53932 451046 53984 451052
rect 53944 266694 53972 451046
rect 54036 353802 54064 451250
rect 55404 422816 55456 422822
rect 55404 422758 55456 422764
rect 55416 412634 55444 422758
rect 55324 412606 55444 412634
rect 55324 410009 55352 412606
rect 55310 410000 55366 410009
rect 55508 409970 55536 604454
rect 66180 576230 66208 616694
rect 71240 616418 71268 619520
rect 77312 616826 77340 619520
rect 77300 616820 77352 616826
rect 77300 616762 77352 616768
rect 78496 616820 78548 616826
rect 78496 616762 78548 616768
rect 71228 616412 71280 616418
rect 71228 616354 71280 616360
rect 78508 604110 78536 616762
rect 80440 616758 80468 619520
rect 80428 616752 80480 616758
rect 80428 616694 80480 616700
rect 81348 616752 81400 616758
rect 81348 616694 81400 616700
rect 78588 616072 78640 616078
rect 78588 616014 78640 616020
rect 78496 604104 78548 604110
rect 78496 604046 78548 604052
rect 66168 576224 66220 576230
rect 66168 576166 66220 576172
rect 78600 566234 78628 616014
rect 79232 599072 79284 599078
rect 79232 599014 79284 599020
rect 78588 566228 78640 566234
rect 78588 566170 78640 566176
rect 75918 566128 75974 566137
rect 75918 566063 75974 566072
rect 75932 565962 75960 566063
rect 75920 565956 75972 565962
rect 75920 565898 75972 565904
rect 76288 565956 76340 565962
rect 76288 565898 76340 565904
rect 59452 539436 59504 539442
rect 59452 539378 59504 539384
rect 59176 539232 59228 539238
rect 59176 539174 59228 539180
rect 59188 507890 59216 539174
rect 59176 507884 59228 507890
rect 59176 507826 59228 507832
rect 55310 409935 55312 409944
rect 55364 409935 55366 409944
rect 55496 409964 55548 409970
rect 55312 409906 55364 409912
rect 55496 409906 55548 409912
rect 54024 353796 54076 353802
rect 54024 353738 54076 353744
rect 53932 266688 53984 266694
rect 53932 266630 53984 266636
rect 53840 222692 53892 222698
rect 53840 222634 53892 222640
rect 54668 222692 54720 222698
rect 54668 222634 54720 222640
rect 54680 220017 54708 222634
rect 55034 220552 55090 220561
rect 55034 220487 55036 220496
rect 55088 220487 55090 220496
rect 55036 220458 55088 220464
rect 54666 220008 54722 220017
rect 54722 219966 54970 219994
rect 54666 219943 54722 219952
rect 54680 219883 54708 219943
rect 53748 219496 53800 219502
rect 53748 219438 53800 219444
rect 55508 219366 55536 409906
rect 57164 409426 57376 409442
rect 57152 409420 57388 409426
rect 57204 409414 57336 409420
rect 57152 409362 57204 409368
rect 57336 409362 57388 409368
rect 56876 409352 56928 409358
rect 56876 409294 56928 409300
rect 56692 409216 56744 409222
rect 56692 409158 56744 409164
rect 56704 356658 56732 409158
rect 56888 409018 56916 409294
rect 56876 409012 56928 409018
rect 56876 408954 56928 408960
rect 56692 356652 56744 356658
rect 56692 356594 56744 356600
rect 59464 237522 59492 539378
rect 59636 539232 59688 539238
rect 59636 539174 59688 539180
rect 59648 287910 59676 539174
rect 75932 524754 75960 565898
rect 76300 565865 76328 565898
rect 76286 565856 76342 565865
rect 76286 565791 76342 565800
rect 75920 524748 75972 524754
rect 75920 524690 75972 524696
rect 64788 447840 64840 447846
rect 64788 447782 64840 447788
rect 64800 313274 64828 447782
rect 67364 422884 67416 422890
rect 67364 422826 67416 422832
rect 67376 400654 67404 422826
rect 67088 400648 67140 400654
rect 67364 400648 67416 400654
rect 67088 400590 67140 400596
rect 67362 400616 67364 400625
rect 67456 400648 67508 400654
rect 67416 400616 67418 400625
rect 67100 356046 67128 400590
rect 67640 400648 67692 400654
rect 67456 400590 67508 400596
rect 67546 400616 67602 400625
rect 67362 400551 67418 400560
rect 67468 364334 67496 400590
rect 67602 400596 67640 400602
rect 67602 400590 67692 400596
rect 67602 400574 67680 400590
rect 67546 400551 67602 400560
rect 67640 400512 67692 400518
rect 67640 400454 67692 400460
rect 67652 400353 67680 400454
rect 67638 400344 67694 400353
rect 67638 400279 67694 400288
rect 71872 378888 71924 378894
rect 71872 378830 71924 378836
rect 70584 378752 70636 378758
rect 70584 378694 70636 378700
rect 67468 364306 67588 364334
rect 67088 356040 67140 356046
rect 67088 355982 67140 355988
rect 67560 355910 67588 364306
rect 67548 355904 67600 355910
rect 67548 355846 67600 355852
rect 67560 355366 67588 355846
rect 67548 355360 67600 355366
rect 67548 355302 67600 355308
rect 64788 313268 64840 313274
rect 64788 313210 64840 313216
rect 61108 304904 61160 304910
rect 61108 304846 61160 304852
rect 59636 287904 59688 287910
rect 59636 287846 59688 287852
rect 59452 237516 59504 237522
rect 59452 237458 59504 237464
rect 61120 236366 61148 304846
rect 70596 292466 70624 378694
rect 71884 306066 71912 378830
rect 71872 306060 71924 306066
rect 71872 306002 71924 306008
rect 70584 292460 70636 292466
rect 70584 292402 70636 292408
rect 78128 264172 78180 264178
rect 78128 264114 78180 264120
rect 77852 264104 77904 264110
rect 77852 264046 77904 264052
rect 77864 236706 77892 264046
rect 77852 236700 77904 236706
rect 77852 236642 77904 236648
rect 77864 236366 77892 236642
rect 61108 236360 61160 236366
rect 61108 236302 61160 236308
rect 77852 236360 77904 236366
rect 77852 236302 77904 236308
rect 61476 236292 61528 236298
rect 61476 236234 61528 236240
rect 61488 236065 61516 236234
rect 62488 236224 62540 236230
rect 62486 236192 62488 236201
rect 62540 236192 62542 236201
rect 62486 236127 62542 236136
rect 61474 236056 61530 236065
rect 61474 235991 61530 236000
rect 61844 223168 61896 223174
rect 61844 223110 61896 223116
rect 61856 222329 61884 223110
rect 68560 222420 68612 222426
rect 68560 222362 68612 222368
rect 61842 222320 61898 222329
rect 61842 222255 61898 222264
rect 61856 219994 61884 222255
rect 68282 220008 68338 220017
rect 61594 219966 61884 219994
rect 68218 219966 68282 219994
rect 68572 219994 68600 222362
rect 75182 222320 75238 222329
rect 75182 222255 75238 222264
rect 75196 219994 75224 222255
rect 77760 220448 77812 220454
rect 77760 220390 77812 220396
rect 68338 219966 68600 219994
rect 74842 219966 75224 219994
rect 68282 219943 68338 219952
rect 68296 219883 68324 219943
rect 77772 219745 77800 220390
rect 77758 219736 77814 219745
rect 77758 219671 77814 219680
rect 78140 219366 78168 264114
rect 79244 263974 79272 599014
rect 81360 528358 81388 616694
rect 83384 616010 83412 619520
rect 83372 616004 83424 616010
rect 83372 615946 83424 615952
rect 86512 615494 86540 619520
rect 92400 616865 92428 619520
rect 92386 616856 92442 616865
rect 92386 616791 92442 616800
rect 95528 615942 95556 619520
rect 95516 615936 95568 615942
rect 95516 615878 95568 615884
rect 98472 615874 98500 619520
rect 101600 616622 101628 619520
rect 101588 616616 101640 616622
rect 101588 616558 101640 616564
rect 104544 616214 104572 619520
rect 106740 616684 106792 616690
rect 106740 616626 106792 616632
rect 103520 616208 103572 616214
rect 103520 616150 103572 616156
rect 104532 616208 104584 616214
rect 104532 616150 104584 616156
rect 98460 615868 98512 615874
rect 98460 615810 98512 615816
rect 86512 615466 86908 615494
rect 82728 557184 82780 557190
rect 82728 557126 82780 557132
rect 81348 528352 81400 528358
rect 81348 528294 81400 528300
rect 79784 339176 79836 339182
rect 79784 339118 79836 339124
rect 79232 263968 79284 263974
rect 79232 263910 79284 263916
rect 79796 220794 79824 339118
rect 82740 222834 82768 557126
rect 86880 265810 86908 615466
rect 101404 558952 101456 558958
rect 101404 558894 101456 558900
rect 93768 493196 93820 493202
rect 93768 493138 93820 493144
rect 93780 473686 93808 493138
rect 93768 473680 93820 473686
rect 93768 473622 93820 473628
rect 93768 473544 93820 473550
rect 93766 473512 93768 473521
rect 97080 473544 97132 473550
rect 93820 473512 93822 473521
rect 97080 473486 97132 473492
rect 93766 473447 93822 473456
rect 93308 473408 93360 473414
rect 93308 473350 93360 473356
rect 93676 473408 93728 473414
rect 93676 473350 93728 473356
rect 88340 446752 88392 446758
rect 88340 446694 88392 446700
rect 88352 359378 88380 446694
rect 91468 434308 91520 434314
rect 91468 434250 91520 434256
rect 91480 433401 91508 434250
rect 91466 433392 91522 433401
rect 91466 433327 91522 433336
rect 91480 425134 91508 433327
rect 91468 425128 91520 425134
rect 91468 425070 91520 425076
rect 92388 425128 92440 425134
rect 92388 425070 92440 425076
rect 89260 423360 89312 423366
rect 89260 423302 89312 423308
rect 89272 384402 89300 423302
rect 92400 423026 92428 425070
rect 92388 423020 92440 423026
rect 92388 422962 92440 422968
rect 89444 409896 89496 409902
rect 89444 409838 89496 409844
rect 89456 384538 89484 409838
rect 92296 409284 92348 409290
rect 92296 409226 92348 409232
rect 90640 409216 90692 409222
rect 90640 409158 90692 409164
rect 89444 384532 89496 384538
rect 89444 384474 89496 384480
rect 89260 384396 89312 384402
rect 89260 384338 89312 384344
rect 88800 384260 88852 384266
rect 88800 384202 88852 384208
rect 88812 384033 88840 384202
rect 89076 384192 89128 384198
rect 89076 384134 89128 384140
rect 89168 384192 89220 384198
rect 89168 384134 89220 384140
rect 88798 384024 88854 384033
rect 88798 383959 88854 383968
rect 88340 359372 88392 359378
rect 88340 359314 88392 359320
rect 89088 334150 89116 384134
rect 89076 334144 89128 334150
rect 89076 334086 89128 334092
rect 89180 273766 89208 384134
rect 89260 381064 89312 381070
rect 89260 381006 89312 381012
rect 89272 356726 89300 381006
rect 90652 356794 90680 409158
rect 90640 356788 90692 356794
rect 90640 356730 90692 356736
rect 89260 356720 89312 356726
rect 89260 356662 89312 356668
rect 89272 356590 89300 356662
rect 89260 356584 89312 356590
rect 90652 356561 90680 356730
rect 89260 356526 89312 356532
rect 90638 356552 90694 356561
rect 90638 356487 90694 356496
rect 89168 273760 89220 273766
rect 89168 273702 89220 273708
rect 92308 270298 92336 409226
rect 93320 326194 93348 473350
rect 93492 359304 93544 359310
rect 93492 359246 93544 359252
rect 93504 326194 93532 359246
rect 93308 326188 93360 326194
rect 93308 326130 93360 326136
rect 93492 326188 93544 326194
rect 93492 326130 93544 326136
rect 92938 288144 92994 288153
rect 92938 288079 92940 288088
rect 92992 288079 92994 288088
rect 93122 288144 93178 288153
rect 93122 288079 93124 288088
rect 92940 288050 92992 288056
rect 93176 288079 93178 288088
rect 93124 288050 93176 288056
rect 92296 270292 92348 270298
rect 92296 270234 92348 270240
rect 92308 269958 92336 270234
rect 92296 269952 92348 269958
rect 92296 269894 92348 269900
rect 86868 265804 86920 265810
rect 86868 265746 86920 265752
rect 93688 223106 93716 473350
rect 95884 425128 95936 425134
rect 95884 425070 95936 425076
rect 95608 415200 95660 415206
rect 95608 415142 95660 415148
rect 95620 374746 95648 415142
rect 95792 378820 95844 378826
rect 95792 378762 95844 378768
rect 95608 374740 95660 374746
rect 95608 374682 95660 374688
rect 95804 374542 95832 378762
rect 95792 374536 95844 374542
rect 95792 374478 95844 374484
rect 95896 229094 95924 425070
rect 95976 384804 96028 384810
rect 95976 384746 96028 384752
rect 95988 374610 96016 384746
rect 95976 374604 96028 374610
rect 95976 374546 96028 374552
rect 95896 229066 96108 229094
rect 93676 223100 93728 223106
rect 93676 223042 93728 223048
rect 95056 222896 95108 222902
rect 95056 222838 95108 222844
rect 81808 222828 81860 222834
rect 81808 222770 81860 222776
rect 82728 222828 82780 222834
rect 82728 222770 82780 222776
rect 79784 220788 79836 220794
rect 79784 220730 79836 220736
rect 79322 220688 79378 220697
rect 79322 220623 79378 220632
rect 79416 220652 79468 220658
rect 79336 220590 79364 220623
rect 79416 220594 79468 220600
rect 79324 220584 79376 220590
rect 79324 220526 79376 220532
rect 79428 220017 79456 220594
rect 79414 220008 79470 220017
rect 81820 219994 81848 222770
rect 81466 219966 81848 219994
rect 94502 220008 94558 220017
rect 79414 219943 79470 219952
rect 95068 219994 95096 222838
rect 94558 219966 95096 219994
rect 94502 219943 94558 219952
rect 96080 219570 96108 229066
rect 97092 220794 97120 473486
rect 99656 411052 99708 411058
rect 99656 410994 99708 411000
rect 99840 411052 99892 411058
rect 99840 410994 99892 411000
rect 99668 348498 99696 410994
rect 99852 410582 99880 410994
rect 99840 410576 99892 410582
rect 99840 410518 99892 410524
rect 99852 349110 99880 410518
rect 99840 349104 99892 349110
rect 99840 349046 99892 349052
rect 100668 349104 100720 349110
rect 100720 349052 100800 349058
rect 100668 349046 100800 349052
rect 99852 348566 99880 349046
rect 100680 349030 100800 349046
rect 99840 348560 99892 348566
rect 99840 348502 99892 348508
rect 99656 348492 99708 348498
rect 99656 348434 99708 348440
rect 100772 345014 100800 349030
rect 100944 348288 100996 348294
rect 100944 348230 100996 348236
rect 100772 344986 100892 345014
rect 98736 263968 98788 263974
rect 98736 263910 98788 263916
rect 98748 263673 98776 263910
rect 98734 263664 98790 263673
rect 98734 263599 98790 263608
rect 100864 224602 100892 344986
rect 100852 224596 100904 224602
rect 100852 224538 100904 224544
rect 100956 224505 100984 348230
rect 100942 224496 100998 224505
rect 100942 224431 100998 224440
rect 100956 224398 100984 224431
rect 100944 224392 100996 224398
rect 100944 224334 100996 224340
rect 101416 222630 101444 558894
rect 101496 415472 101548 415478
rect 101496 415414 101548 415420
rect 101404 222624 101456 222630
rect 101404 222566 101456 222572
rect 97080 220788 97132 220794
rect 97080 220730 97132 220736
rect 96620 220584 96672 220590
rect 96620 220526 96672 220532
rect 96068 219564 96120 219570
rect 96068 219506 96120 219512
rect 96632 219473 96660 220526
rect 101416 220017 101444 222566
rect 101402 220008 101458 220017
rect 101338 219966 101402 219994
rect 101402 219943 101458 219952
rect 101416 219883 101444 219943
rect 87786 219464 87842 219473
rect 96618 219464 96674 219473
rect 87842 219422 88090 219450
rect 87786 219399 87842 219408
rect 96618 219399 96674 219408
rect 101508 219366 101536 415414
rect 103532 384198 103560 616150
rect 106752 584730 106780 616626
rect 110616 616350 110644 619520
rect 113744 616826 113772 619520
rect 113732 616820 113784 616826
rect 113732 616762 113784 616768
rect 114376 616820 114428 616826
rect 114376 616762 114428 616768
rect 114100 616752 114152 616758
rect 114100 616694 114152 616700
rect 110604 616344 110656 616350
rect 110604 616286 110656 616292
rect 111892 590980 111944 590986
rect 111892 590922 111944 590928
rect 106740 584724 106792 584730
rect 106740 584666 106792 584672
rect 111904 467226 111932 590922
rect 112536 527468 112588 527474
rect 112536 527410 112588 527416
rect 112444 473612 112496 473618
rect 112444 473554 112496 473560
rect 111892 467220 111944 467226
rect 111892 467162 111944 467168
rect 112350 446992 112406 447001
rect 112260 446956 112312 446962
rect 112350 446927 112352 446936
rect 112260 446898 112312 446904
rect 112404 446927 112406 446936
rect 112352 446898 112404 446904
rect 108304 384736 108356 384742
rect 108304 384678 108356 384684
rect 103520 384192 103572 384198
rect 103518 384160 103520 384169
rect 103572 384160 103574 384169
rect 103518 384095 103574 384104
rect 106372 356652 106424 356658
rect 106372 356594 106424 356600
rect 106188 353320 106240 353326
rect 106188 353262 106240 353268
rect 106200 336122 106228 353262
rect 106188 336116 106240 336122
rect 106188 336058 106240 336064
rect 106384 335986 106412 356594
rect 106372 335980 106424 335986
rect 106372 335922 106424 335928
rect 108316 286958 108344 384678
rect 112168 295724 112220 295730
rect 112168 295666 112220 295672
rect 112180 295633 112208 295666
rect 112166 295624 112222 295633
rect 112166 295559 112222 295568
rect 108304 286952 108356 286958
rect 108304 286894 108356 286900
rect 103426 266928 103482 266937
rect 103426 266863 103482 266872
rect 103440 248441 103468 266863
rect 103426 248432 103482 248441
rect 103426 248367 103482 248376
rect 103426 238640 103482 238649
rect 103426 238575 103482 238584
rect 103440 229129 103468 238575
rect 103426 229120 103482 229129
rect 103426 229055 103482 229064
rect 103426 228984 103482 228993
rect 103426 228919 103482 228928
rect 103440 224913 103468 228919
rect 103426 224904 103482 224913
rect 103426 224839 103482 224848
rect 112272 223038 112300 446898
rect 112456 446894 112484 473554
rect 112444 446888 112496 446894
rect 112444 446830 112496 446836
rect 112548 410650 112576 527410
rect 113088 524544 113140 524550
rect 113088 524486 113140 524492
rect 112996 467424 113048 467430
rect 112996 467366 113048 467372
rect 113008 467090 113036 467366
rect 112996 467084 113048 467090
rect 112996 467026 113048 467032
rect 112628 467016 112680 467022
rect 112628 466958 112680 466964
rect 112640 443494 112668 466958
rect 112812 466948 112864 466954
rect 112812 466890 112864 466896
rect 112628 443488 112680 443494
rect 112628 443430 112680 443436
rect 112536 410644 112588 410650
rect 112536 410586 112588 410592
rect 112824 410553 112852 466890
rect 113008 410650 113036 467026
rect 112996 410644 113048 410650
rect 112996 410586 113048 410592
rect 112810 410544 112866 410553
rect 112810 410479 112866 410488
rect 112824 410446 112852 410479
rect 112812 410440 112864 410446
rect 112812 410382 112864 410388
rect 112824 410310 112852 410382
rect 112812 410304 112864 410310
rect 112812 410246 112864 410252
rect 112536 295724 112588 295730
rect 112536 295666 112588 295672
rect 112260 223032 112312 223038
rect 112260 222974 112312 222980
rect 112548 220726 112576 295666
rect 112536 220720 112588 220726
rect 112536 220662 112588 220668
rect 107660 220652 107712 220658
rect 107660 220594 107712 220600
rect 107672 219994 107700 220594
rect 107672 219966 107962 219994
rect 113008 219366 113036 410586
rect 113100 410514 113128 524486
rect 113088 410508 113140 410514
rect 113088 410450 113140 410456
rect 114112 405618 114140 616694
rect 114100 405612 114152 405618
rect 114100 405554 114152 405560
rect 114388 219366 114416 616762
rect 115952 335374 115980 619534
rect 116504 619426 116532 619534
rect 116646 619520 116758 620960
rect 119774 619520 119886 620960
rect 122718 619520 122830 620960
rect 125846 619520 125958 620960
rect 128790 619520 128902 620960
rect 131734 619520 131846 620960
rect 134862 619520 134974 620960
rect 137806 619520 137918 620960
rect 140934 619520 141046 620960
rect 143878 619520 143990 620960
rect 147006 619520 147118 620960
rect 149950 619520 150062 620960
rect 153078 619520 153190 620960
rect 156022 619520 156134 620960
rect 159150 619520 159262 620960
rect 162094 619520 162206 620960
rect 165222 619520 165334 620960
rect 168166 619520 168278 620960
rect 171110 619520 171222 620960
rect 174238 619520 174350 620960
rect 177182 619520 177294 620960
rect 180310 619520 180422 620960
rect 183254 619520 183366 620960
rect 186382 619520 186494 620960
rect 189326 619520 189438 620960
rect 192454 619520 192566 620960
rect 194612 619534 195284 619562
rect 116688 619426 116716 619520
rect 116504 619398 116716 619426
rect 119816 615494 119844 619520
rect 122760 616282 122788 619520
rect 125888 616690 125916 619520
rect 125876 616684 125928 616690
rect 125876 616626 125928 616632
rect 128832 616486 128860 619520
rect 131776 616690 131804 619520
rect 134524 616888 134576 616894
rect 134524 616830 134576 616836
rect 131764 616684 131816 616690
rect 131764 616626 131816 616632
rect 128820 616480 128872 616486
rect 128820 616422 128872 616428
rect 122748 616276 122800 616282
rect 122748 616218 122800 616224
rect 119816 615466 120028 615494
rect 120000 547874 120028 615466
rect 121368 578944 121420 578950
rect 121368 578886 121420 578892
rect 119908 547846 120028 547874
rect 119528 547460 119580 547466
rect 119528 547402 119580 547408
rect 119540 541754 119568 547402
rect 119528 541748 119580 541754
rect 119528 541690 119580 541696
rect 119908 538214 119936 547846
rect 120080 541544 120132 541550
rect 119986 541512 120042 541521
rect 120080 541486 120132 541492
rect 119986 541447 119988 541456
rect 120040 541447 120042 541456
rect 119988 541418 120040 541424
rect 119908 538186 120028 538214
rect 119620 414792 119672 414798
rect 119620 414734 119672 414740
rect 119632 414089 119660 414734
rect 119618 414080 119674 414089
rect 119618 414015 119674 414024
rect 120000 401742 120028 538186
rect 120092 465254 120120 541486
rect 121000 526176 121052 526182
rect 121000 526118 121052 526124
rect 120080 465248 120132 465254
rect 120080 465190 120132 465196
rect 121012 422958 121040 526118
rect 121000 422952 121052 422958
rect 121000 422894 121052 422900
rect 119988 401736 120040 401742
rect 119988 401678 120040 401684
rect 115940 335368 115992 335374
rect 115940 335310 115992 335316
rect 117780 326188 117832 326194
rect 117780 326130 117832 326136
rect 114468 295724 114520 295730
rect 114468 295666 114520 295672
rect 114480 295633 114508 295666
rect 114466 295624 114522 295633
rect 114466 295559 114522 295568
rect 117596 256352 117648 256358
rect 117596 256294 117648 256300
rect 117608 252890 117636 256294
rect 117596 252884 117648 252890
rect 117596 252826 117648 252832
rect 117792 252686 117820 326130
rect 117780 252680 117832 252686
rect 117780 252622 117832 252628
rect 121380 219994 121408 578886
rect 123392 561604 123444 561610
rect 123392 561546 123444 561552
rect 121828 546848 121880 546854
rect 121828 546790 121880 546796
rect 121840 528562 121868 546790
rect 123300 541680 123352 541686
rect 123298 541648 123300 541657
rect 123352 541648 123354 541657
rect 123298 541583 123354 541592
rect 121828 528556 121880 528562
rect 121828 528498 121880 528504
rect 123404 220794 123432 561546
rect 133696 429548 133748 429554
rect 133696 429490 133748 429496
rect 133708 423502 133736 429490
rect 132592 423496 132644 423502
rect 132592 423438 132644 423444
rect 133696 423496 133748 423502
rect 133696 423438 133748 423444
rect 133880 423496 133932 423502
rect 133880 423438 133932 423444
rect 133972 423496 134024 423502
rect 133972 423438 134024 423444
rect 134156 423496 134208 423502
rect 134156 423438 134208 423444
rect 132604 384334 132632 423438
rect 133892 422618 133920 423438
rect 133984 423162 134012 423438
rect 133972 423156 134024 423162
rect 133972 423098 134024 423104
rect 134168 423094 134196 423438
rect 134340 423360 134392 423366
rect 134340 423302 134392 423308
rect 134156 423088 134208 423094
rect 134156 423030 134208 423036
rect 133880 422612 133932 422618
rect 133880 422554 133932 422560
rect 132592 384328 132644 384334
rect 132590 384296 132592 384305
rect 132644 384296 132646 384305
rect 132590 384231 132646 384240
rect 132408 384192 132460 384198
rect 132408 384134 132460 384140
rect 130384 383240 130436 383246
rect 130384 383182 130436 383188
rect 125876 273964 125928 273970
rect 125876 273906 125928 273912
rect 125784 261248 125836 261254
rect 125322 261216 125378 261225
rect 125784 261190 125836 261196
rect 125322 261151 125378 261160
rect 125336 260914 125364 261151
rect 125796 260914 125824 261190
rect 125888 261050 125916 273906
rect 125876 261044 125928 261050
rect 125876 260986 125928 260992
rect 125874 260944 125930 260953
rect 125324 260908 125376 260914
rect 125324 260850 125376 260856
rect 125784 260908 125836 260914
rect 125874 260879 125876 260888
rect 125784 260850 125836 260856
rect 125928 260879 125930 260888
rect 125876 260850 125928 260856
rect 123392 220788 123444 220794
rect 123392 220730 123444 220736
rect 123404 220697 123432 220730
rect 123390 220688 123446 220697
rect 123390 220623 123446 220632
rect 125336 220250 125364 260850
rect 125796 220522 125824 260850
rect 126980 230784 127032 230790
rect 126980 230726 127032 230732
rect 126992 223582 127020 230726
rect 126980 223576 127032 223582
rect 126980 223518 127032 223524
rect 127532 223576 127584 223582
rect 127532 223518 127584 223524
rect 125784 220516 125836 220522
rect 125784 220458 125836 220464
rect 125324 220244 125376 220250
rect 125324 220186 125376 220192
rect 121210 219966 121408 219994
rect 127544 219994 127572 223518
rect 127544 219966 127834 219994
rect 114926 219464 114982 219473
rect 114586 219422 114926 219450
rect 130396 219434 130424 383182
rect 132420 296002 132448 384134
rect 131120 295996 131172 296002
rect 131120 295938 131172 295944
rect 132408 295996 132460 296002
rect 132408 295938 132460 295944
rect 131132 295798 131160 295938
rect 131120 295792 131172 295798
rect 131120 295734 131172 295740
rect 134352 283762 134380 423302
rect 134340 283756 134392 283762
rect 134340 283698 134392 283704
rect 130476 261316 130528 261322
rect 130476 261258 130528 261264
rect 130488 261225 130516 261258
rect 130474 261216 130530 261225
rect 130474 261151 130530 261160
rect 131578 260944 131634 260953
rect 131578 260879 131580 260888
rect 131632 260879 131634 260888
rect 131580 260850 131632 260856
rect 133236 236700 133288 236706
rect 133236 236642 133288 236648
rect 133248 220590 133276 236642
rect 134536 223514 134564 616830
rect 134904 616554 134932 619520
rect 137848 616554 137876 619520
rect 143920 616826 143948 619520
rect 143908 616820 143960 616826
rect 143908 616762 143960 616768
rect 134892 616548 134944 616554
rect 134892 616490 134944 616496
rect 137836 616548 137888 616554
rect 137836 616490 137888 616496
rect 153844 616480 153896 616486
rect 153844 616422 153896 616428
rect 136548 616276 136600 616282
rect 136548 616218 136600 616224
rect 136560 417178 136588 616218
rect 153200 615868 153252 615874
rect 153200 615810 153252 615816
rect 143816 615800 143868 615806
rect 143816 615742 143868 615748
rect 137192 613896 137244 613902
rect 137192 613838 137244 613844
rect 136548 417172 136600 417178
rect 136548 417114 136600 417120
rect 136548 381540 136600 381546
rect 136548 381482 136600 381488
rect 136560 380934 136588 381482
rect 136088 380928 136140 380934
rect 136088 380870 136140 380876
rect 136548 380928 136600 380934
rect 136548 380870 136600 380876
rect 135904 280288 135956 280294
rect 135904 280230 135956 280236
rect 135916 227186 135944 280230
rect 136100 229094 136128 380870
rect 136008 229066 136128 229094
rect 136008 227186 136036 229066
rect 137204 227730 137232 613838
rect 142436 600704 142488 600710
rect 142436 600646 142488 600652
rect 142068 584044 142120 584050
rect 142068 583986 142120 583992
rect 140780 446888 140832 446894
rect 140780 446830 140832 446836
rect 137928 335912 137980 335918
rect 137928 335854 137980 335860
rect 137940 292398 137968 335854
rect 140792 307154 140820 446830
rect 140780 307148 140832 307154
rect 140780 307090 140832 307096
rect 140778 307048 140834 307057
rect 140778 306983 140780 306992
rect 140832 306983 140834 306992
rect 140780 306954 140832 306960
rect 140872 306944 140924 306950
rect 140872 306886 140924 306892
rect 141240 306944 141292 306950
rect 141240 306886 141292 306892
rect 137928 292392 137980 292398
rect 137928 292334 137980 292340
rect 137192 227724 137244 227730
rect 137192 227666 137244 227672
rect 137192 227588 137244 227594
rect 137192 227530 137244 227536
rect 135628 227180 135680 227186
rect 135628 227122 135680 227128
rect 135904 227180 135956 227186
rect 135904 227122 135956 227128
rect 135996 227180 136048 227186
rect 135996 227122 136048 227128
rect 135640 227089 135668 227122
rect 137204 227118 137232 227530
rect 136548 227112 136600 227118
rect 135626 227080 135682 227089
rect 135626 227015 135682 227024
rect 136546 227080 136548 227089
rect 137192 227112 137244 227118
rect 136600 227080 136602 227089
rect 137192 227054 137244 227060
rect 136546 227015 136602 227024
rect 137204 226681 137232 227054
rect 137190 226672 137246 226681
rect 137190 226607 137246 226616
rect 134524 223508 134576 223514
rect 134524 223450 134576 223456
rect 133236 220584 133288 220590
rect 133236 220526 133288 220532
rect 134536 220017 134564 223450
rect 137940 220522 137968 292334
rect 140884 222834 140912 306886
rect 141252 267918 141280 306886
rect 141240 267912 141292 267918
rect 141240 267854 141292 267860
rect 142080 223582 142108 583986
rect 142344 448588 142396 448594
rect 142344 448530 142396 448536
rect 142356 429418 142384 448530
rect 142448 429554 142476 600646
rect 143080 434920 143132 434926
rect 143080 434862 143132 434868
rect 142436 429548 142488 429554
rect 142436 429490 142488 429496
rect 142344 429412 142396 429418
rect 142344 429354 142396 429360
rect 142448 384402 142476 429490
rect 142436 384396 142488 384402
rect 142436 384338 142488 384344
rect 143092 365430 143120 434862
rect 143828 412826 143856 615742
rect 152372 443692 152424 443698
rect 152372 443634 152424 443640
rect 152280 443148 152332 443154
rect 152280 443090 152332 443096
rect 152292 441614 152320 443090
rect 152384 443057 152412 443634
rect 152464 443624 152516 443630
rect 152464 443566 152516 443572
rect 152370 443048 152426 443057
rect 152370 442983 152426 442992
rect 152292 441586 152412 441614
rect 143816 412820 143868 412826
rect 143816 412762 143868 412768
rect 152384 374542 152412 441586
rect 152476 415546 152504 443566
rect 153016 443012 153068 443018
rect 153016 442954 153068 442960
rect 152464 415540 152516 415546
rect 152464 415482 152516 415488
rect 152372 374536 152424 374542
rect 152372 374478 152424 374484
rect 143080 365424 143132 365430
rect 143078 365392 143080 365401
rect 143132 365392 143134 365401
rect 143078 365327 143134 365336
rect 143092 365158 143120 365327
rect 143080 365152 143132 365158
rect 143080 365094 143132 365100
rect 153028 362642 153056 442954
rect 153016 362636 153068 362642
rect 153016 362578 153068 362584
rect 141424 223576 141476 223582
rect 141424 223518 141476 223524
rect 142068 223576 142120 223582
rect 142068 223518 142120 223524
rect 140872 222828 140924 222834
rect 140872 222770 140924 222776
rect 137928 220516 137980 220522
rect 137928 220458 137980 220464
rect 134522 220008 134578 220017
rect 134458 219966 134522 219994
rect 141436 219994 141464 223518
rect 147772 223100 147824 223106
rect 147772 223042 147824 223048
rect 147784 219994 147812 223042
rect 153212 222698 153240 615810
rect 153476 525088 153528 525094
rect 153476 525030 153528 525036
rect 153384 304768 153436 304774
rect 153384 304710 153436 304716
rect 153396 229838 153424 304710
rect 153488 229838 153516 525030
rect 153856 502246 153884 616422
rect 156064 605834 156092 619520
rect 162136 616078 162164 619520
rect 177224 616321 177252 619520
rect 183296 616486 183324 619520
rect 183284 616480 183336 616486
rect 183284 616422 183336 616428
rect 184572 616480 184624 616486
rect 184572 616422 184624 616428
rect 177210 616312 177266 616321
rect 177210 616247 177266 616256
rect 162124 616072 162176 616078
rect 162124 616014 162176 616020
rect 160744 616004 160796 616010
rect 160744 615946 160796 615952
rect 155972 605806 156092 605834
rect 153844 502240 153896 502246
rect 153844 502182 153896 502188
rect 155972 236230 156000 605806
rect 158904 599208 158956 599214
rect 158904 599150 158956 599156
rect 158444 565888 158496 565894
rect 158444 565830 158496 565836
rect 157430 543824 157486 543833
rect 157248 543788 157300 543794
rect 157430 543759 157432 543768
rect 157248 543730 157300 543736
rect 157484 543759 157486 543768
rect 157524 543788 157576 543794
rect 157432 543730 157484 543736
rect 157524 543730 157576 543736
rect 157260 514214 157288 543730
rect 157536 524618 157564 543730
rect 158456 540530 158484 565830
rect 158444 540524 158496 540530
rect 158444 540466 158496 540472
rect 158628 540524 158680 540530
rect 158628 540466 158680 540472
rect 158640 540326 158668 540466
rect 158720 540388 158772 540394
rect 158720 540330 158772 540336
rect 158812 540388 158864 540394
rect 158812 540330 158864 540336
rect 158628 540320 158680 540326
rect 158628 540262 158680 540268
rect 158640 524822 158668 540262
rect 158732 526182 158760 540330
rect 158720 526176 158772 526182
rect 158720 526118 158772 526124
rect 158628 524816 158680 524822
rect 158628 524758 158680 524764
rect 157524 524612 157576 524618
rect 157524 524554 157576 524560
rect 157248 514208 157300 514214
rect 157248 514150 157300 514156
rect 158824 261322 158852 540330
rect 158916 273970 158944 599150
rect 158996 599140 159048 599146
rect 158996 599082 159048 599088
rect 158904 273964 158956 273970
rect 158904 273906 158956 273912
rect 159008 273902 159036 599082
rect 159088 540388 159140 540394
rect 159088 540330 159140 540336
rect 159100 539617 159128 540330
rect 159086 539608 159142 539617
rect 159086 539543 159142 539552
rect 159088 434240 159140 434246
rect 159088 434182 159140 434188
rect 159100 273970 159128 434182
rect 159088 273964 159140 273970
rect 159088 273906 159140 273912
rect 159272 273964 159324 273970
rect 159272 273906 159324 273912
rect 158996 273896 159048 273902
rect 159284 273873 159312 273906
rect 158996 273838 159048 273844
rect 159270 273864 159326 273873
rect 158812 261316 158864 261322
rect 158812 261258 158864 261264
rect 155960 236224 156012 236230
rect 155960 236166 156012 236172
rect 153384 229832 153436 229838
rect 153476 229832 153528 229838
rect 153384 229774 153436 229780
rect 153474 229800 153476 229809
rect 153528 229800 153530 229809
rect 153474 229735 153530 229744
rect 159008 229094 159036 273838
rect 159270 273799 159326 273808
rect 159008 229066 159128 229094
rect 153200 222692 153252 222698
rect 153200 222634 153252 222640
rect 154028 222692 154080 222698
rect 154028 222634 154080 222640
rect 154040 220017 154068 222634
rect 159100 220726 159128 229066
rect 159088 220720 159140 220726
rect 159088 220662 159140 220668
rect 159100 220289 159128 220662
rect 159086 220280 159142 220289
rect 159086 220215 159142 220224
rect 141082 219966 141464 219994
rect 147706 219966 147812 219994
rect 154026 220008 154082 220017
rect 134522 219943 134578 219952
rect 160756 219994 160784 615946
rect 167736 615936 167788 615942
rect 167736 615878 167788 615884
rect 167276 613896 167328 613902
rect 167276 613838 167328 613844
rect 167644 613896 167696 613902
rect 167644 613838 167696 613844
rect 167288 483818 167316 613838
rect 167276 483812 167328 483818
rect 167276 483754 167328 483760
rect 167458 228304 167514 228313
rect 167458 228239 167460 228248
rect 167512 228239 167514 228248
rect 167460 228210 167512 228216
rect 167184 228200 167236 228206
rect 167368 228200 167420 228206
rect 167184 228142 167236 228148
rect 167366 228168 167368 228177
rect 167420 228168 167422 228177
rect 162768 220584 162820 220590
rect 162768 220526 162820 220532
rect 154082 219966 154330 219994
rect 160756 219980 160954 219994
rect 160756 219966 160968 219980
rect 154026 219943 154082 219952
rect 134536 219883 134564 219943
rect 154040 219883 154068 219943
rect 160940 219450 160968 219966
rect 162780 219706 162808 220526
rect 167196 219978 167224 228142
rect 167366 228103 167422 228112
rect 167656 227730 167684 613838
rect 167644 227724 167696 227730
rect 167644 227666 167696 227672
rect 167656 227118 167684 227666
rect 167644 227112 167696 227118
rect 167644 227054 167696 227060
rect 167748 219994 167776 615878
rect 175740 613964 175792 613970
rect 175740 613906 175792 613912
rect 175648 613828 175700 613834
rect 175648 613770 175700 613776
rect 167920 613760 167972 613766
rect 167920 613702 167972 613708
rect 167932 469810 167960 613702
rect 167920 469804 167972 469810
rect 167920 469746 167972 469752
rect 170404 460964 170456 460970
rect 170404 460906 170456 460912
rect 170416 402966 170444 460906
rect 175660 448458 175688 613770
rect 175752 448526 175780 613906
rect 182088 612808 182140 612814
rect 182088 612750 182140 612756
rect 180432 578740 180484 578746
rect 180432 578682 180484 578688
rect 176936 536852 176988 536858
rect 176936 536794 176988 536800
rect 175740 448520 175792 448526
rect 175740 448462 175792 448468
rect 176016 448520 176068 448526
rect 176016 448462 176068 448468
rect 175556 448452 175608 448458
rect 175556 448394 175608 448400
rect 175648 448452 175700 448458
rect 175648 448394 175700 448400
rect 170404 402960 170456 402966
rect 170404 402902 170456 402908
rect 167828 393780 167880 393786
rect 167828 393722 167880 393728
rect 167840 228410 167868 393722
rect 175568 333198 175596 448394
rect 175556 333192 175608 333198
rect 175556 333134 175608 333140
rect 167828 228404 167880 228410
rect 167828 228346 167880 228352
rect 175660 227254 175688 448394
rect 175752 332858 175780 448462
rect 176028 333130 176056 448462
rect 176016 333124 176068 333130
rect 176016 333066 176068 333072
rect 175740 332852 175792 332858
rect 175740 332794 175792 332800
rect 176948 277914 176976 536794
rect 177028 513732 177080 513738
rect 177028 513674 177080 513680
rect 177040 383994 177068 513674
rect 178316 448452 178368 448458
rect 178316 448394 178368 448400
rect 177304 409352 177356 409358
rect 177304 409294 177356 409300
rect 177028 383988 177080 383994
rect 177028 383930 177080 383936
rect 177210 383888 177266 383897
rect 177316 383858 177344 409294
rect 177210 383823 177212 383832
rect 177264 383823 177266 383832
rect 177304 383852 177356 383858
rect 177212 383794 177264 383800
rect 177304 383794 177356 383800
rect 176936 277908 176988 277914
rect 176936 277850 176988 277856
rect 175832 228200 175884 228206
rect 175830 228168 175832 228177
rect 175884 228168 175886 228177
rect 175830 228103 175886 228112
rect 175648 227248 175700 227254
rect 175648 227190 175700 227196
rect 178328 220658 178356 448394
rect 180444 362642 180472 578682
rect 180432 362636 180484 362642
rect 180432 362578 180484 362584
rect 180062 362536 180118 362545
rect 180062 362471 180064 362480
rect 180116 362471 180118 362480
rect 180064 362442 180116 362448
rect 182100 317422 182128 612750
rect 184584 601458 184612 616422
rect 184572 601452 184624 601458
rect 184572 601394 184624 601400
rect 190368 500064 190420 500070
rect 190368 500006 190420 500012
rect 190380 499633 190408 500006
rect 190366 499624 190422 499633
rect 190366 499559 190422 499568
rect 194612 475386 194640 619534
rect 195256 619426 195284 619534
rect 195398 619520 195510 620960
rect 198526 619520 198638 620960
rect 201470 619520 201582 620960
rect 204598 619520 204710 620960
rect 207542 619520 207654 620960
rect 210486 619520 210598 620960
rect 213614 619520 213726 620960
rect 216558 619520 216670 620960
rect 219686 619520 219798 620960
rect 222630 619520 222742 620960
rect 225758 619520 225870 620960
rect 228702 619520 228814 620960
rect 231830 619520 231942 620960
rect 234774 619520 234886 620960
rect 237902 619520 238014 620960
rect 240846 619520 240958 620960
rect 243974 619520 244086 620960
rect 246918 619520 247030 620960
rect 249862 619520 249974 620960
rect 252990 619520 253102 620960
rect 255934 619520 256046 620960
rect 259062 619520 259174 620960
rect 262006 619520 262118 620960
rect 265134 619520 265246 620960
rect 267752 619534 267964 619562
rect 195440 619426 195468 619520
rect 195256 619398 195468 619426
rect 198568 615806 198596 619520
rect 210528 615806 210556 619520
rect 198556 615800 198608 615806
rect 198556 615742 198608 615748
rect 210516 615800 210568 615806
rect 210516 615742 210568 615748
rect 211068 615800 211120 615806
rect 211068 615742 211120 615748
rect 196440 600840 196492 600846
rect 196440 600782 196492 600788
rect 196452 572082 196480 600782
rect 206008 596556 206060 596562
rect 206008 596498 206060 596504
rect 205454 596456 205510 596465
rect 205454 596391 205510 596400
rect 205468 596358 205496 596391
rect 205456 596352 205508 596358
rect 205456 596294 205508 596300
rect 205824 596352 205876 596358
rect 205916 596352 205968 596358
rect 205824 596294 205876 596300
rect 205914 596320 205916 596329
rect 205968 596320 205970 596329
rect 203984 587104 204036 587110
rect 203984 587046 204036 587052
rect 201500 583976 201552 583982
rect 201500 583918 201552 583924
rect 201512 583817 201540 583918
rect 201960 583840 202012 583846
rect 201498 583808 201554 583817
rect 201960 583782 202012 583788
rect 201498 583743 201554 583752
rect 196440 572076 196492 572082
rect 196440 572018 196492 572024
rect 194600 475380 194652 475386
rect 194600 475322 194652 475328
rect 198280 471300 198332 471306
rect 198280 471242 198332 471248
rect 198464 471300 198516 471306
rect 198464 471242 198516 471248
rect 194784 470960 194836 470966
rect 194784 470902 194836 470908
rect 194796 467226 194824 470902
rect 198292 470665 198320 471242
rect 198278 470656 198334 470665
rect 198278 470591 198334 470600
rect 194784 467220 194836 467226
rect 194784 467162 194836 467168
rect 195060 466948 195112 466954
rect 195060 466890 195112 466896
rect 184572 428256 184624 428262
rect 184572 428198 184624 428204
rect 182088 317416 182140 317422
rect 182088 317358 182140 317364
rect 184584 316034 184612 428198
rect 193680 354272 193732 354278
rect 193680 354214 193732 354220
rect 193692 353394 193720 354214
rect 194600 353456 194652 353462
rect 194598 353424 194600 353433
rect 194652 353424 194654 353433
rect 193588 353388 193640 353394
rect 193588 353330 193640 353336
rect 193680 353388 193732 353394
rect 194598 353359 194654 353368
rect 193680 353330 193732 353336
rect 193600 335782 193628 353330
rect 193864 353320 193916 353326
rect 193864 353262 193916 353268
rect 193588 335776 193640 335782
rect 193588 335718 193640 335724
rect 184492 316006 184612 316034
rect 184492 312118 184520 316006
rect 184480 312112 184532 312118
rect 184480 312054 184532 312060
rect 180800 307148 180852 307154
rect 180800 307090 180852 307096
rect 180812 259282 180840 307090
rect 193876 300966 193904 353262
rect 193864 300960 193916 300966
rect 193864 300902 193916 300908
rect 195072 291242 195100 466890
rect 195244 439748 195296 439754
rect 195244 439690 195296 439696
rect 195256 354414 195284 439690
rect 198476 409970 198504 471242
rect 198464 409964 198516 409970
rect 198464 409906 198516 409912
rect 200488 384260 200540 384266
rect 200488 384202 200540 384208
rect 199660 383852 199712 383858
rect 199660 383794 199712 383800
rect 199672 383654 199700 383794
rect 199752 383784 199804 383790
rect 199752 383726 199804 383732
rect 200120 383784 200172 383790
rect 200500 383738 200528 384202
rect 200172 383732 200528 383738
rect 200120 383726 200528 383732
rect 199660 383648 199712 383654
rect 199660 383590 199712 383596
rect 199764 376754 199792 383726
rect 200132 383710 200528 383726
rect 199764 376726 199976 376754
rect 195244 354408 195296 354414
rect 195244 354350 195296 354356
rect 195428 354408 195480 354414
rect 195428 354350 195480 354356
rect 195440 353394 195468 354350
rect 195428 353388 195480 353394
rect 195428 353330 195480 353336
rect 195060 291236 195112 291242
rect 195060 291178 195112 291184
rect 180800 259276 180852 259282
rect 180800 259218 180852 259224
rect 180984 259276 181036 259282
rect 180984 259218 181036 259224
rect 180890 259176 180946 259185
rect 180890 259111 180892 259120
rect 180944 259111 180946 259120
rect 180892 259082 180944 259088
rect 180800 259072 180852 259078
rect 180800 259014 180852 259020
rect 180812 258641 180840 259014
rect 180798 258632 180854 258641
rect 180798 258567 180854 258576
rect 180996 238754 181024 259218
rect 181260 259072 181312 259078
rect 181260 259014 181312 259020
rect 181272 257582 181300 259014
rect 181260 257576 181312 257582
rect 181260 257518 181312 257524
rect 180812 238726 181024 238754
rect 180812 228206 180840 238726
rect 180800 228200 180852 228206
rect 180800 228142 180852 228148
rect 187608 223304 187660 223310
rect 187608 223246 187660 223252
rect 178316 220652 178368 220658
rect 178316 220594 178368 220600
rect 167184 219972 167236 219978
rect 167578 219966 167776 219994
rect 167184 219914 167236 219920
rect 162768 219700 162820 219706
rect 162768 219642 162820 219648
rect 162780 219609 162808 219642
rect 162766 219600 162822 219609
rect 162766 219535 162822 219544
rect 161294 219464 161350 219473
rect 160940 219436 161294 219450
rect 114926 219399 114982 219408
rect 130384 219428 130436 219434
rect 160954 219422 161294 219436
rect 167748 219450 167776 219966
rect 187146 220008 187202 220017
rect 187620 219994 187648 223246
rect 194416 223236 194468 223242
rect 194416 223178 194468 223184
rect 187202 219966 187648 219994
rect 193770 220008 193826 220017
rect 187146 219943 187202 219952
rect 194428 219994 194456 223178
rect 199948 222766 199976 376726
rect 201972 301102 202000 583782
rect 203996 559162 204024 587046
rect 203984 559156 204036 559162
rect 203984 559098 204036 559104
rect 204352 558952 204404 558958
rect 204352 558894 204404 558900
rect 203064 473408 203116 473414
rect 203064 473350 203116 473356
rect 203076 417450 203104 473350
rect 203064 417444 203116 417450
rect 203064 417386 203116 417392
rect 201960 301096 202012 301102
rect 201960 301038 202012 301044
rect 204364 230858 204392 558894
rect 205272 423156 205324 423162
rect 205272 423098 205324 423104
rect 204996 296200 205048 296206
rect 204996 296142 205048 296148
rect 204352 230852 204404 230858
rect 204352 230794 204404 230800
rect 200396 223032 200448 223038
rect 200396 222974 200448 222980
rect 199936 222760 199988 222766
rect 199936 222702 199988 222708
rect 193826 219966 194456 219994
rect 200408 219994 200436 222974
rect 205008 220794 205036 296142
rect 204996 220788 205048 220794
rect 204996 220730 205048 220736
rect 205008 220658 205036 220730
rect 205284 220658 205312 423098
rect 205364 423088 205416 423094
rect 205364 423030 205416 423036
rect 205376 220946 205404 423030
rect 205640 413636 205692 413642
rect 205640 413578 205692 413584
rect 205376 220918 205588 220946
rect 204996 220652 205048 220658
rect 204996 220594 205048 220600
rect 205180 220652 205232 220658
rect 205180 220594 205232 220600
rect 205272 220652 205324 220658
rect 205272 220594 205324 220600
rect 200408 219966 200698 219994
rect 193770 219943 193826 219952
rect 205192 219638 205220 220594
rect 205284 220454 205312 220594
rect 205376 220590 205404 220918
rect 205456 220788 205508 220794
rect 205456 220730 205508 220736
rect 205364 220584 205416 220590
rect 205364 220526 205416 220532
rect 205468 220538 205496 220730
rect 205560 220674 205588 220918
rect 205652 220794 205680 413578
rect 205836 222698 205864 596294
rect 205914 596255 205970 596264
rect 206020 584458 206048 596498
rect 206008 584452 206060 584458
rect 206008 584394 206060 584400
rect 206020 583914 206048 584394
rect 206008 583908 206060 583914
rect 206008 583850 206060 583856
rect 208308 565956 208360 565962
rect 208308 565898 208360 565904
rect 208320 498166 208348 565898
rect 208308 498160 208360 498166
rect 208308 498102 208360 498108
rect 208582 498128 208638 498137
rect 208320 497894 208348 498102
rect 208582 498063 208584 498072
rect 208636 498063 208638 498072
rect 208584 498034 208636 498040
rect 208308 497888 208360 497894
rect 208308 497830 208360 497836
rect 208492 492040 208544 492046
rect 208492 491982 208544 491988
rect 207112 491904 207164 491910
rect 207112 491846 207164 491852
rect 207020 355360 207072 355366
rect 207020 355302 207072 355308
rect 207032 262478 207060 355302
rect 207124 273222 207152 491846
rect 208504 467226 208532 491982
rect 208492 467220 208544 467226
rect 208492 467162 208544 467168
rect 207204 465452 207256 465458
rect 207204 465394 207256 465400
rect 207112 273216 207164 273222
rect 207112 273158 207164 273164
rect 207216 262614 207244 465394
rect 211080 397526 211108 615742
rect 213656 615494 213684 619520
rect 222672 616078 222700 619520
rect 222660 616072 222712 616078
rect 222660 616014 222712 616020
rect 216220 615868 216272 615874
rect 216220 615810 216272 615816
rect 213656 615466 213868 615494
rect 213840 571946 213868 615466
rect 213828 571940 213880 571946
rect 213828 571882 213880 571888
rect 211068 397520 211120 397526
rect 211068 397462 211120 397468
rect 214564 389224 214616 389230
rect 214564 389166 214616 389172
rect 207204 262608 207256 262614
rect 207204 262550 207256 262556
rect 207020 262472 207072 262478
rect 207388 262472 207440 262478
rect 207020 262414 207072 262420
rect 207386 262440 207388 262449
rect 207440 262440 207442 262449
rect 207386 262375 207442 262384
rect 214576 229094 214604 389166
rect 214748 370184 214800 370190
rect 214748 370126 214800 370132
rect 214760 369889 214788 370126
rect 214746 369880 214802 369889
rect 214746 369815 214802 369824
rect 216232 231538 216260 615810
rect 228744 615494 228772 619520
rect 231872 616865 231900 619520
rect 234816 616865 234844 619520
rect 240888 616865 240916 619520
rect 231858 616856 231914 616865
rect 231858 616791 231914 616800
rect 234802 616856 234858 616865
rect 234802 616791 234858 616800
rect 240874 616856 240930 616865
rect 240874 616791 240930 616800
rect 233424 616072 233476 616078
rect 233424 616014 233476 616020
rect 228744 615466 229048 615494
rect 228456 606892 228508 606898
rect 228456 606834 228508 606840
rect 228468 606121 228496 606834
rect 228454 606112 228510 606121
rect 228454 606047 228510 606056
rect 221464 540456 221516 540462
rect 221464 540398 221516 540404
rect 220544 355904 220596 355910
rect 220544 355846 220596 355852
rect 218702 337648 218758 337657
rect 218702 337583 218758 337592
rect 218716 337550 218744 337583
rect 218704 337544 218756 337550
rect 218704 337486 218756 337492
rect 218520 337408 218572 337414
rect 218520 337350 218572 337356
rect 216220 231532 216272 231538
rect 216220 231474 216272 231480
rect 214392 229066 214604 229094
rect 207388 223440 207440 223446
rect 207388 223382 207440 223388
rect 205824 222692 205876 222698
rect 205824 222634 205876 222640
rect 207400 222329 207428 223382
rect 214392 222465 214420 229066
rect 214378 222456 214434 222465
rect 214378 222391 214434 222400
rect 207386 222320 207442 222329
rect 207386 222255 207442 222264
rect 205640 220788 205692 220794
rect 205640 220730 205692 220736
rect 205732 220788 205784 220794
rect 205732 220730 205784 220736
rect 205744 220674 205772 220730
rect 205560 220646 205772 220674
rect 205468 220522 205588 220538
rect 205468 220516 205600 220522
rect 205468 220510 205548 220516
rect 205548 220458 205600 220464
rect 205272 220448 205324 220454
rect 205272 220390 205324 220396
rect 207400 219994 207428 222255
rect 209042 220824 209098 220833
rect 209042 220759 209044 220768
rect 209096 220759 209098 220768
rect 209044 220730 209096 220736
rect 213184 220448 213236 220454
rect 213182 220416 213184 220425
rect 213236 220416 213238 220425
rect 213182 220351 213238 220360
rect 214392 219994 214420 222391
rect 207322 219966 207428 219994
rect 213946 219966 214420 219994
rect 205180 219632 205232 219638
rect 205178 219600 205180 219609
rect 205232 219600 205234 219609
rect 205178 219535 205234 219544
rect 167918 219464 167974 219473
rect 167748 219422 167918 219450
rect 161294 219399 161350 219408
rect 167918 219399 167974 219408
rect 173990 219464 174046 219473
rect 181166 219464 181222 219473
rect 174046 219422 174202 219450
rect 180826 219422 181166 219450
rect 173990 219399 174046 219408
rect 181166 219399 181222 219408
rect 130384 219370 130436 219376
rect 218532 219366 218560 337350
rect 220556 254930 220584 355846
rect 221476 271182 221504 540398
rect 229020 537742 229048 615466
rect 231860 606484 231912 606490
rect 231860 606426 231912 606432
rect 231872 572150 231900 606426
rect 233436 600302 233464 616014
rect 247592 615800 247644 615806
rect 247592 615742 247644 615748
rect 237840 611584 237892 611590
rect 237840 611526 237892 611532
rect 236460 607368 236512 607374
rect 236460 607310 236512 607316
rect 233424 600296 233476 600302
rect 233424 600238 233476 600244
rect 233332 576904 233384 576910
rect 233332 576846 233384 576852
rect 231860 572144 231912 572150
rect 231860 572086 231912 572092
rect 231872 548690 231900 572086
rect 231860 548684 231912 548690
rect 231860 548626 231912 548632
rect 232136 548548 232188 548554
rect 232136 548490 232188 548496
rect 229008 537736 229060 537742
rect 229008 537678 229060 537684
rect 228916 473544 228968 473550
rect 228916 473486 228968 473492
rect 224408 465384 224460 465390
rect 224408 465326 224460 465332
rect 224420 443630 224448 465326
rect 224408 443624 224460 443630
rect 224408 443566 224460 443572
rect 227904 281580 227956 281586
rect 227904 281522 227956 281528
rect 221464 271176 221516 271182
rect 221464 271118 221516 271124
rect 220544 254924 220596 254930
rect 220544 254866 220596 254872
rect 219806 254824 219862 254833
rect 219806 254759 219808 254768
rect 219860 254759 219862 254768
rect 219808 254730 219860 254736
rect 219256 254720 219308 254726
rect 219254 254688 219256 254697
rect 219308 254688 219310 254697
rect 219254 254623 219310 254632
rect 227916 248414 227944 281522
rect 228928 267918 228956 473486
rect 232148 415274 232176 548490
rect 232136 415268 232188 415274
rect 232136 415210 232188 415216
rect 232688 384260 232740 384266
rect 232688 384202 232740 384208
rect 232320 348356 232372 348362
rect 232320 348298 232372 348304
rect 231032 337476 231084 337482
rect 231032 337418 231084 337424
rect 231044 337385 231072 337418
rect 231030 337376 231086 337385
rect 231030 337311 231086 337320
rect 228916 267912 228968 267918
rect 228916 267854 228968 267860
rect 229098 267880 229154 267889
rect 229098 267815 229154 267824
rect 229112 267782 229140 267815
rect 229100 267776 229152 267782
rect 229100 267718 229152 267724
rect 232332 250986 232360 348298
rect 232700 344146 232728 384202
rect 233344 344282 233372 576846
rect 236472 571130 236500 607310
rect 236460 571124 236512 571130
rect 236460 571066 236512 571072
rect 236472 570790 236500 571066
rect 237852 570994 237880 611526
rect 247604 596698 247632 615742
rect 259104 615641 259132 619520
rect 262048 615942 262076 619520
rect 265176 616758 265204 619520
rect 265164 616752 265216 616758
rect 265164 616694 265216 616700
rect 262036 615936 262088 615942
rect 262036 615878 262088 615884
rect 259090 615632 259146 615641
rect 259090 615567 259146 615576
rect 263876 607232 263928 607238
rect 263876 607174 263928 607180
rect 247592 596692 247644 596698
rect 247592 596634 247644 596640
rect 262496 584452 262548 584458
rect 262496 584394 262548 584400
rect 247684 576972 247736 576978
rect 247684 576914 247736 576920
rect 237564 570988 237616 570994
rect 237564 570930 237616 570936
rect 237840 570988 237892 570994
rect 237840 570930 237892 570936
rect 236460 570784 236512 570790
rect 236460 570726 236512 570732
rect 237576 567194 237604 570930
rect 237576 567166 237696 567194
rect 233700 566024 233752 566030
rect 233700 565966 233752 565972
rect 233712 371890 233740 565966
rect 233792 498092 233844 498098
rect 233792 498034 233844 498040
rect 233700 371884 233752 371890
rect 233700 371826 233752 371832
rect 233712 371793 233740 371826
rect 233698 371784 233754 371793
rect 233698 371719 233754 371728
rect 233804 371686 233832 498034
rect 237380 492040 237432 492046
rect 237380 491982 237432 491988
rect 237392 489870 237420 491982
rect 237380 489864 237432 489870
rect 237380 489806 237432 489812
rect 237668 487286 237696 567166
rect 244924 518560 244976 518566
rect 244924 518502 244976 518508
rect 238208 489864 238260 489870
rect 238208 489806 238260 489812
rect 237656 487280 237708 487286
rect 237656 487222 237708 487228
rect 238220 480146 238248 489806
rect 238208 480140 238260 480146
rect 238208 480082 238260 480088
rect 238484 480004 238536 480010
rect 238484 479946 238536 479952
rect 233792 371680 233844 371686
rect 233792 371622 233844 371628
rect 233332 344276 233384 344282
rect 233332 344218 233384 344224
rect 232688 344140 232740 344146
rect 232688 344082 232740 344088
rect 232700 259282 232728 344082
rect 232964 343936 233016 343942
rect 232964 343878 233016 343884
rect 232688 259276 232740 259282
rect 232688 259218 232740 259224
rect 232320 250980 232372 250986
rect 232320 250922 232372 250928
rect 227916 248386 228128 248414
rect 228100 223582 228128 248386
rect 228088 223576 228140 223582
rect 228088 223518 228140 223524
rect 227536 222352 227588 222358
rect 227536 222294 227588 222300
rect 226982 220008 227038 220017
rect 227548 219994 227576 222294
rect 227038 219966 227576 219994
rect 226982 219943 227038 219952
rect 232976 219366 233004 343878
rect 235264 220652 235316 220658
rect 235264 220594 235316 220600
rect 235276 220017 235304 220594
rect 238496 220114 238524 479946
rect 239036 424584 239088 424590
rect 239036 424526 239088 424532
rect 239048 223378 239076 424526
rect 244464 423428 244516 423434
rect 244464 423370 244516 423376
rect 244372 360392 244424 360398
rect 244372 360334 244424 360340
rect 243084 311976 243136 311982
rect 243084 311918 243136 311924
rect 240140 292256 240192 292262
rect 240140 292198 240192 292204
rect 239036 223372 239088 223378
rect 239036 223314 239088 223320
rect 240152 222601 240180 292198
rect 243096 283694 243124 311918
rect 244384 295322 244412 360334
rect 244372 295316 244424 295322
rect 244372 295258 244424 295264
rect 244476 283898 244504 423370
rect 244464 283892 244516 283898
rect 244464 283834 244516 283840
rect 243084 283688 243136 283694
rect 243084 283630 243136 283636
rect 244476 283558 244504 283834
rect 244464 283552 244516 283558
rect 244464 283494 244516 283500
rect 240322 232520 240378 232529
rect 240322 232455 240324 232464
rect 240376 232455 240378 232464
rect 240324 232426 240376 232432
rect 240138 222592 240194 222601
rect 240138 222527 240194 222536
rect 238484 220108 238536 220114
rect 238484 220050 238536 220056
rect 235262 220008 235318 220017
rect 235262 219943 235318 219952
rect 240152 219994 240180 222527
rect 240152 219966 240442 219994
rect 240152 219745 240180 219966
rect 240138 219736 240194 219745
rect 240138 219671 240194 219680
rect 234158 219464 234214 219473
rect 233818 219422 234158 219450
rect 234158 219399 234214 219408
rect 20536 219360 20588 219366
rect 20536 219302 20588 219308
rect 21548 219360 21600 219366
rect 21548 219302 21600 219308
rect 22928 219360 22980 219366
rect 22928 219302 22980 219308
rect 55496 219360 55548 219366
rect 55496 219302 55548 219308
rect 78128 219360 78180 219366
rect 78128 219302 78180 219308
rect 101496 219360 101548 219366
rect 101496 219302 101548 219308
rect 112996 219360 113048 219366
rect 112996 219302 113048 219308
rect 114376 219360 114428 219366
rect 114376 219302 114428 219308
rect 218520 219360 218572 219366
rect 232964 219360 233016 219366
rect 218520 219302 218572 219308
rect 220266 219328 220322 219337
rect 220322 219286 220570 219314
rect 244936 219337 244964 518502
rect 247696 507482 247724 576914
rect 258908 561672 258960 561678
rect 258908 561614 258960 561620
rect 255688 559020 255740 559026
rect 255688 558962 255740 558968
rect 247684 507476 247736 507482
rect 247684 507418 247736 507424
rect 247592 507272 247644 507278
rect 247592 507214 247644 507220
rect 247604 467430 247632 507214
rect 248144 507136 248196 507142
rect 248144 507078 248196 507084
rect 247592 467424 247644 467430
rect 247592 467366 247644 467372
rect 248156 364682 248184 507078
rect 255596 496392 255648 496398
rect 255596 496334 255648 496340
rect 255608 495854 255636 496334
rect 255700 495922 255728 558962
rect 255688 495916 255740 495922
rect 255688 495858 255740 495864
rect 255596 495848 255648 495854
rect 255596 495790 255648 495796
rect 248328 489796 248380 489802
rect 248328 489738 248380 489744
rect 248144 364676 248196 364682
rect 248144 364618 248196 364624
rect 248236 273964 248288 273970
rect 248236 273906 248288 273912
rect 248248 273873 248276 273906
rect 248234 273864 248290 273873
rect 248234 273799 248290 273808
rect 247132 222828 247184 222834
rect 247132 222770 247184 222776
rect 247144 219994 247172 222770
rect 247066 219966 247172 219994
rect 248340 219366 248368 489738
rect 249432 489728 249484 489734
rect 249432 489670 249484 489676
rect 248696 276140 248748 276146
rect 248696 276082 248748 276088
rect 248604 276072 248656 276078
rect 248604 276014 248656 276020
rect 248616 273902 248644 276014
rect 248604 273896 248656 273902
rect 248604 273838 248656 273844
rect 248708 220726 248736 276082
rect 248696 220720 248748 220726
rect 248696 220662 248748 220668
rect 249444 219366 249472 489670
rect 255608 465322 255636 495790
rect 255596 465316 255648 465322
rect 255596 465258 255648 465264
rect 254216 457224 254268 457230
rect 254216 457166 254268 457172
rect 254124 457088 254176 457094
rect 254124 457030 254176 457036
rect 254136 412690 254164 457030
rect 254124 412684 254176 412690
rect 254124 412626 254176 412632
rect 254136 410990 254164 412626
rect 254124 410984 254176 410990
rect 254124 410926 254176 410932
rect 253112 410372 253164 410378
rect 253112 410314 253164 410320
rect 253124 399430 253152 410314
rect 253112 399424 253164 399430
rect 253112 399366 253164 399372
rect 252560 267776 252612 267782
rect 252560 267718 252612 267724
rect 252572 222562 252600 267718
rect 254228 250918 254256 457166
rect 255700 288114 255728 495858
rect 257068 415336 257120 415342
rect 257068 415278 257120 415284
rect 257080 344146 257108 415278
rect 258920 413914 258948 561614
rect 260656 548616 260708 548622
rect 260656 548558 260708 548564
rect 260668 513874 260696 548558
rect 262508 525230 262536 584394
rect 262770 525328 262826 525337
rect 262770 525263 262772 525272
rect 262824 525263 262826 525272
rect 262772 525234 262824 525240
rect 262496 525224 262548 525230
rect 262680 525224 262732 525230
rect 262496 525166 262548 525172
rect 262678 525192 262680 525201
rect 262732 525192 262734 525201
rect 260656 513868 260708 513874
rect 260656 513810 260708 513816
rect 259184 513664 259236 513670
rect 259184 513606 259236 513612
rect 258908 413908 258960 413914
rect 258908 413850 258960 413856
rect 257436 412684 257488 412690
rect 257436 412626 257488 412632
rect 257068 344140 257120 344146
rect 257068 344082 257120 344088
rect 255688 288108 255740 288114
rect 255688 288050 255740 288056
rect 257160 283552 257212 283558
rect 257160 283494 257212 283500
rect 254216 250912 254268 250918
rect 254216 250854 254268 250860
rect 255962 223272 256018 223281
rect 255962 223207 255964 223216
rect 256016 223207 256018 223216
rect 255964 223178 256016 223184
rect 252560 222556 252612 222562
rect 252560 222498 252612 222504
rect 253388 222556 253440 222562
rect 253388 222498 253440 222504
rect 249708 220720 249760 220726
rect 249708 220662 249760 220668
rect 249720 219774 249748 220662
rect 253400 220017 253428 222498
rect 257172 220590 257200 283494
rect 257252 250912 257304 250918
rect 257252 250854 257304 250860
rect 257264 220590 257292 250854
rect 257448 220658 257476 412626
rect 258920 220726 258948 413850
rect 259196 383994 259224 513606
rect 259368 479936 259420 479942
rect 259368 479878 259420 479884
rect 259380 478922 259408 479878
rect 259368 478916 259420 478922
rect 259368 478858 259420 478864
rect 259380 470594 259408 478858
rect 259288 470566 259408 470594
rect 259184 383988 259236 383994
rect 259184 383930 259236 383936
rect 259092 295860 259144 295866
rect 259092 295802 259144 295808
rect 258908 220720 258960 220726
rect 258908 220662 258960 220668
rect 259104 220658 259132 295802
rect 259184 222420 259236 222426
rect 259184 222362 259236 222368
rect 259196 220697 259224 222362
rect 259288 220726 259316 470566
rect 262508 415342 262536 525166
rect 262678 525127 262734 525136
rect 263692 485580 263744 485586
rect 263692 485522 263744 485528
rect 263704 485382 263732 485522
rect 263888 485518 263916 607174
rect 265072 545148 265124 545154
rect 265072 545090 265124 545096
rect 264060 485648 264112 485654
rect 264060 485590 264112 485596
rect 263876 485512 263928 485518
rect 263876 485454 263928 485460
rect 264072 485466 264100 485590
rect 263508 485376 263560 485382
rect 263508 485318 263560 485324
rect 263692 485376 263744 485382
rect 263692 485318 263744 485324
rect 263784 485376 263836 485382
rect 263784 485318 263836 485324
rect 263520 471374 263548 485318
rect 263508 471368 263560 471374
rect 263508 471310 263560 471316
rect 263704 436121 263732 485318
rect 263690 436112 263746 436121
rect 263690 436047 263746 436056
rect 263704 434858 263732 436047
rect 263692 434852 263744 434858
rect 263692 434794 263744 434800
rect 262496 415336 262548 415342
rect 262496 415278 262548 415284
rect 259552 378888 259604 378894
rect 259552 378830 259604 378836
rect 259460 295588 259512 295594
rect 259460 295530 259512 295536
rect 259276 220720 259328 220726
rect 259182 220688 259238 220697
rect 257436 220652 257488 220658
rect 257436 220594 257488 220600
rect 259092 220652 259144 220658
rect 259276 220662 259328 220668
rect 259472 220658 259500 295530
rect 259564 229094 259592 378830
rect 263600 301640 263652 301646
rect 263600 301582 263652 301588
rect 261116 301504 261168 301510
rect 261116 301446 261168 301452
rect 262312 301504 262364 301510
rect 262312 301446 262364 301452
rect 261128 300937 261156 301446
rect 261114 300928 261170 300937
rect 261114 300863 261170 300872
rect 262324 296070 262352 301446
rect 262312 296064 262364 296070
rect 262312 296006 262364 296012
rect 263612 283762 263640 301582
rect 263600 283756 263652 283762
rect 263600 283698 263652 283704
rect 263612 279410 263640 283698
rect 263600 279404 263652 279410
rect 263600 279346 263652 279352
rect 263796 255270 263824 485318
rect 263888 365430 263916 485454
rect 264072 485450 264192 485466
rect 264072 485444 264204 485450
rect 264072 485438 264152 485444
rect 263876 365424 263928 365430
rect 263876 365366 263928 365372
rect 264072 365362 264100 485438
rect 264152 485386 264204 485392
rect 264060 365356 264112 365362
rect 264060 365298 264112 365304
rect 264612 308576 264664 308582
rect 264612 308518 264664 308524
rect 264624 279478 264652 308518
rect 264612 279472 264664 279478
rect 264612 279414 264664 279420
rect 263784 255264 263836 255270
rect 263784 255206 263836 255212
rect 263796 254726 263824 255206
rect 263784 254720 263836 254726
rect 263784 254662 263836 254668
rect 260656 252612 260708 252618
rect 260656 252554 260708 252560
rect 260668 229094 260696 252554
rect 259564 229066 259684 229094
rect 260668 229066 260788 229094
rect 259656 220658 259684 229066
rect 260760 224954 260788 229066
rect 260668 224926 260788 224954
rect 260668 223530 260696 224926
rect 260840 223576 260892 223582
rect 260668 223524 260840 223530
rect 260668 223518 260892 223524
rect 260668 223502 260880 223518
rect 260472 223304 260524 223310
rect 260472 223246 260524 223252
rect 260564 223304 260616 223310
rect 260564 223246 260616 223252
rect 260484 222578 260512 223246
rect 260576 223174 260604 223246
rect 260668 223174 260696 223502
rect 260746 223272 260802 223281
rect 260746 223207 260748 223216
rect 260800 223207 260802 223216
rect 260748 223178 260800 223184
rect 260564 223168 260616 223174
rect 260564 223110 260616 223116
rect 260656 223168 260708 223174
rect 260656 223110 260708 223116
rect 260484 222550 260788 222578
rect 260656 222420 260708 222426
rect 260656 222362 260708 222368
rect 259182 220623 259184 220632
rect 259092 220594 259144 220600
rect 259236 220623 259238 220632
rect 259460 220652 259512 220658
rect 259184 220594 259236 220600
rect 259460 220594 259512 220600
rect 259644 220652 259696 220658
rect 259644 220594 259696 220600
rect 257160 220584 257212 220590
rect 257160 220526 257212 220532
rect 257252 220584 257304 220590
rect 257252 220526 257304 220532
rect 253386 220008 253442 220017
rect 253442 219966 253690 219994
rect 253386 219943 253442 219952
rect 253400 219883 253428 219943
rect 249708 219768 249760 219774
rect 249708 219710 249760 219716
rect 257172 219570 257200 220526
rect 257356 220522 257660 220538
rect 257344 220516 257672 220522
rect 257396 220510 257620 220516
rect 257344 220458 257396 220464
rect 257620 220458 257672 220464
rect 257712 220448 257764 220454
rect 257712 220390 257764 220396
rect 257724 219881 257752 220390
rect 257710 219872 257766 219881
rect 257710 219807 257766 219816
rect 259104 219706 259132 220594
rect 259196 220563 259224 220594
rect 259472 219910 259500 220594
rect 259656 220114 259684 220594
rect 259644 220108 259696 220114
rect 259644 220050 259696 220056
rect 260668 219994 260696 222362
rect 260314 219966 260696 219994
rect 259460 219904 259512 219910
rect 259460 219846 259512 219852
rect 259092 219700 259144 219706
rect 259092 219642 259144 219648
rect 257160 219564 257212 219570
rect 257160 219506 257212 219512
rect 260760 219366 260788 222550
rect 265084 220454 265112 545090
rect 267648 514344 267700 514350
rect 267648 514286 267700 514292
rect 266360 279404 266412 279410
rect 266360 279346 266412 279352
rect 266372 251122 266400 279346
rect 266360 251116 266412 251122
rect 266360 251058 266412 251064
rect 266372 248414 266400 251058
rect 266372 248386 266492 248414
rect 266464 229094 266492 248386
rect 267660 229094 267688 514286
rect 267752 433430 267780 619534
rect 267936 619426 267964 619534
rect 268078 619520 268190 620960
rect 271206 619520 271318 620960
rect 274150 619520 274262 620960
rect 277278 619520 277390 620960
rect 280222 619520 280334 620960
rect 283350 619520 283462 620960
rect 286294 619520 286406 620960
rect 289238 619520 289350 620960
rect 291212 619534 292252 619562
rect 268120 619426 268148 619520
rect 267936 619398 268148 619426
rect 274192 616185 274220 619520
rect 274178 616176 274234 616185
rect 274178 616111 274234 616120
rect 277320 616078 277348 619520
rect 277308 616072 277360 616078
rect 277308 616014 277360 616020
rect 268384 615732 268436 615738
rect 268384 615674 268436 615680
rect 268292 553580 268344 553586
rect 268292 553522 268344 553528
rect 268304 553489 268332 553522
rect 268290 553480 268346 553489
rect 268290 553415 268346 553424
rect 267740 433424 267792 433430
rect 267740 433366 267792 433372
rect 268396 259214 268424 615674
rect 280264 615602 280292 619520
rect 285312 616752 285364 616758
rect 285312 616694 285364 616700
rect 281356 616072 281408 616078
rect 281356 616014 281408 616020
rect 280252 615596 280304 615602
rect 280252 615538 280304 615544
rect 268568 553580 268620 553586
rect 268568 553522 268620 553528
rect 268752 553580 268804 553586
rect 268752 553522 268804 553528
rect 268844 553580 268896 553586
rect 268844 553522 268896 553528
rect 268580 553489 268608 553522
rect 268566 553480 268622 553489
rect 268566 553415 268622 553424
rect 268764 337414 268792 553522
rect 268856 471306 268884 553522
rect 279240 548548 279292 548554
rect 279240 548490 279292 548496
rect 273904 540320 273956 540326
rect 273904 540262 273956 540268
rect 273628 526380 273680 526386
rect 273628 526322 273680 526328
rect 268844 471300 268896 471306
rect 268844 471242 268896 471248
rect 268752 337408 268804 337414
rect 268752 337350 268804 337356
rect 273640 287065 273668 526322
rect 273916 306374 273944 540262
rect 276940 513868 276992 513874
rect 276940 513810 276992 513816
rect 276952 492250 276980 513810
rect 276940 492244 276992 492250
rect 276940 492186 276992 492192
rect 276952 492114 276980 492186
rect 276940 492108 276992 492114
rect 276940 492050 276992 492056
rect 276952 489870 276980 492050
rect 277308 491972 277360 491978
rect 277308 491914 277360 491920
rect 277320 491706 277348 491914
rect 277308 491700 277360 491706
rect 277308 491642 277360 491648
rect 276940 489864 276992 489870
rect 276940 489806 276992 489812
rect 279252 415410 279280 548490
rect 281368 442610 281396 616014
rect 281448 615596 281500 615602
rect 281448 615538 281500 615544
rect 281356 442604 281408 442610
rect 281356 442546 281408 442552
rect 281460 436966 281488 615538
rect 283012 610632 283064 610638
rect 283012 610574 283064 610580
rect 283024 610230 283052 610574
rect 283288 610564 283340 610570
rect 283288 610506 283340 610512
rect 283380 610564 283432 610570
rect 283380 610506 283432 610512
rect 283012 610224 283064 610230
rect 283012 610166 283064 610172
rect 281448 436960 281500 436966
rect 281448 436902 281500 436908
rect 281356 432200 281408 432206
rect 281356 432142 281408 432148
rect 281630 432168 281686 432177
rect 279240 415404 279292 415410
rect 279240 415346 279292 415352
rect 279608 415336 279660 415342
rect 279608 415278 279660 415284
rect 279620 383926 279648 415278
rect 281368 413710 281396 432142
rect 281630 432103 281632 432112
rect 281684 432103 281686 432112
rect 281632 432074 281684 432080
rect 282736 432064 282788 432070
rect 282734 432032 282736 432041
rect 282788 432032 282790 432041
rect 282734 431967 282790 431976
rect 281356 413704 281408 413710
rect 281356 413646 281408 413652
rect 279608 383920 279660 383926
rect 279608 383862 279660 383868
rect 274454 380488 274510 380497
rect 274454 380423 274456 380432
rect 274508 380423 274510 380432
rect 274456 380394 274508 380400
rect 282276 325032 282328 325038
rect 282274 325000 282276 325009
rect 282328 325000 282330 325009
rect 282274 324935 282330 324944
rect 273916 306346 274036 306374
rect 273626 287056 273682 287065
rect 273626 286991 273628 287000
rect 273680 286991 273682 287000
rect 273812 287020 273864 287026
rect 273628 286962 273680 286968
rect 273812 286962 273864 286968
rect 273640 286931 273668 286962
rect 273824 261050 273852 286962
rect 274008 286890 274036 306346
rect 274732 293344 274784 293350
rect 274732 293286 274784 293292
rect 273996 286884 274048 286890
rect 273996 286826 274048 286832
rect 274008 285705 274036 286826
rect 273994 285696 274050 285705
rect 273994 285631 274050 285640
rect 273812 261044 273864 261050
rect 273812 260986 273864 260992
rect 268384 259208 268436 259214
rect 268384 259150 268436 259156
rect 274744 251190 274772 293286
rect 274732 251184 274784 251190
rect 274732 251126 274784 251132
rect 283024 229094 283052 610166
rect 283300 400586 283328 610506
rect 283392 610065 283420 610506
rect 283378 610056 283434 610065
rect 283378 609991 283434 610000
rect 285324 570994 285352 616694
rect 289280 615874 289308 619520
rect 289268 615868 289320 615874
rect 289268 615810 289320 615816
rect 291212 579086 291240 619534
rect 292224 619426 292252 619534
rect 292366 619520 292478 620960
rect 295310 619520 295422 620960
rect 298438 619520 298550 620960
rect 301382 619520 301494 620960
rect 304510 619520 304622 620960
rect 307454 619520 307566 620960
rect 310582 619520 310694 620960
rect 313526 619520 313638 620960
rect 316052 619534 316540 619562
rect 292408 619426 292436 619520
rect 292224 619398 292436 619426
rect 295352 616865 295380 619520
rect 295338 616856 295394 616865
rect 295338 616791 295394 616800
rect 298480 615806 298508 619520
rect 310624 616826 310652 619520
rect 299204 616820 299256 616826
rect 299204 616762 299256 616768
rect 310612 616820 310664 616826
rect 310612 616762 310664 616768
rect 311808 616820 311860 616826
rect 311808 616762 311860 616768
rect 313372 616820 313424 616826
rect 313372 616762 313424 616768
rect 298468 615800 298520 615806
rect 298468 615742 298520 615748
rect 291200 579080 291252 579086
rect 291200 579022 291252 579028
rect 285312 570988 285364 570994
rect 285312 570930 285364 570936
rect 290832 525224 290884 525230
rect 290832 525166 290884 525172
rect 289820 518696 289872 518702
rect 289818 518664 289820 518673
rect 289872 518664 289874 518673
rect 290844 518634 290872 525166
rect 291106 518800 291162 518809
rect 291106 518735 291108 518744
rect 291160 518735 291162 518744
rect 291108 518706 291160 518712
rect 289818 518599 289874 518608
rect 290832 518628 290884 518634
rect 290832 518570 290884 518576
rect 290280 495848 290332 495854
rect 290280 495790 290332 495796
rect 290004 428392 290056 428398
rect 290004 428334 290056 428340
rect 283288 400580 283340 400586
rect 283288 400522 283340 400528
rect 266464 229066 266676 229094
rect 266084 220720 266136 220726
rect 266084 220662 266136 220668
rect 266096 220538 266124 220662
rect 266648 220590 266676 229066
rect 267384 229066 267688 229094
rect 282932 229066 283052 229094
rect 266636 220584 266688 220590
rect 266096 220510 266584 220538
rect 266636 220526 266688 220532
rect 266556 220454 266584 220510
rect 265072 220448 265124 220454
rect 265072 220390 265124 220396
rect 266544 220448 266596 220454
rect 266544 220390 266596 220396
rect 264978 219872 265034 219881
rect 265084 219842 265112 220390
rect 266648 220386 266676 220526
rect 266636 220380 266688 220386
rect 266636 220322 266688 220328
rect 266648 219881 266676 220322
rect 267384 219994 267412 229066
rect 280528 223032 280580 223038
rect 280528 222974 280580 222980
rect 280540 220017 280568 222974
rect 282932 220658 282960 229066
rect 289820 224800 289872 224806
rect 289820 224742 289872 224748
rect 289832 224466 289860 224742
rect 290016 224602 290044 428334
rect 290292 225010 290320 495790
rect 297640 475720 297692 475726
rect 297640 475662 297692 475668
rect 293684 434308 293736 434314
rect 293684 434250 293736 434256
rect 293696 369102 293724 434250
rect 293684 369096 293736 369102
rect 293684 369038 293736 369044
rect 296076 353864 296128 353870
rect 296076 353806 296128 353812
rect 296088 283354 296116 353806
rect 297652 283762 297680 475662
rect 297640 283756 297692 283762
rect 297640 283698 297692 283704
rect 296904 283688 296956 283694
rect 296904 283630 296956 283636
rect 296076 283348 296128 283354
rect 296076 283290 296128 283296
rect 296720 283144 296772 283150
rect 296720 283086 296772 283092
rect 296732 282810 296760 283086
rect 296916 283082 296944 283630
rect 297652 283218 297680 283698
rect 297640 283212 297692 283218
rect 297640 283154 297692 283160
rect 296904 283076 296956 283082
rect 296904 283018 296956 283024
rect 296720 282804 296772 282810
rect 296720 282746 296772 282752
rect 296916 282674 296944 283018
rect 296076 282668 296128 282674
rect 296076 282610 296128 282616
rect 296904 282668 296956 282674
rect 296904 282610 296956 282616
rect 296088 282538 296116 282610
rect 296076 282532 296128 282538
rect 296076 282474 296128 282480
rect 296088 270094 296116 282474
rect 296076 270088 296128 270094
rect 296076 270030 296128 270036
rect 298836 269952 298888 269958
rect 298836 269894 298888 269900
rect 298848 256494 298876 269894
rect 299216 256562 299244 616762
rect 310796 606688 310848 606694
rect 310796 606630 310848 606636
rect 310612 556776 310664 556782
rect 310612 556718 310664 556724
rect 309692 514412 309744 514418
rect 309692 514354 309744 514360
rect 308312 432200 308364 432206
rect 308312 432142 308364 432148
rect 308324 375698 308352 432142
rect 309704 375834 309732 514354
rect 309692 375828 309744 375834
rect 309692 375770 309744 375776
rect 308312 375692 308364 375698
rect 308312 375634 308364 375640
rect 309704 375494 309732 375770
rect 309692 375488 309744 375494
rect 309692 375430 309744 375436
rect 310624 334422 310652 556718
rect 310612 334416 310664 334422
rect 310612 334358 310664 334364
rect 310624 334286 310652 334358
rect 310808 334286 310836 606630
rect 311164 549296 311216 549302
rect 311164 549238 311216 549244
rect 310612 334280 310664 334286
rect 310612 334222 310664 334228
rect 310796 334280 310848 334286
rect 310796 334222 310848 334228
rect 310704 271176 310756 271182
rect 310704 271118 310756 271124
rect 310244 267912 310296 267918
rect 310244 267854 310296 267860
rect 299388 266756 299440 266762
rect 299388 266698 299440 266704
rect 299400 256698 299428 266698
rect 299388 256692 299440 256698
rect 299388 256634 299440 256640
rect 299204 256556 299256 256562
rect 299204 256498 299256 256504
rect 298836 256488 298888 256494
rect 298836 256430 298888 256436
rect 310060 256012 310112 256018
rect 310060 255954 310112 255960
rect 303160 250028 303212 250034
rect 303160 249970 303212 249976
rect 303172 249937 303200 249970
rect 303158 249928 303214 249937
rect 303158 249863 303214 249872
rect 290280 225004 290332 225010
rect 290280 224946 290332 224952
rect 290004 224596 290056 224602
rect 290004 224538 290056 224544
rect 289820 224460 289872 224466
rect 289820 224402 289872 224408
rect 289636 224256 289688 224262
rect 289636 224198 289688 224204
rect 289648 223689 289676 224198
rect 289634 223680 289690 223689
rect 289634 223615 289690 223624
rect 299756 222760 299808 222766
rect 299756 222702 299808 222708
rect 286508 222692 286560 222698
rect 286508 222634 286560 222640
rect 282920 220652 282972 220658
rect 282920 220594 282972 220600
rect 280526 220008 280582 220017
rect 266938 219966 267412 219994
rect 280186 219966 280526 219994
rect 280526 219943 280582 219952
rect 280540 219883 280568 219943
rect 266634 219872 266690 219881
rect 264978 219807 264980 219816
rect 265032 219807 265034 219816
rect 265072 219836 265124 219842
rect 264980 219778 265032 219784
rect 266634 219807 266690 219816
rect 265072 219778 265124 219784
rect 282932 219706 282960 220594
rect 286520 219994 286548 222634
rect 299768 219994 299796 222702
rect 286520 219966 286810 219994
rect 299768 219966 300058 219994
rect 282920 219700 282972 219706
rect 282920 219642 282972 219648
rect 273258 219464 273314 219473
rect 293222 219464 293278 219473
rect 273314 219422 273562 219450
rect 273258 219399 273314 219408
rect 293278 219422 293434 219450
rect 293222 219399 293278 219408
rect 248328 219360 248380 219366
rect 232964 219302 233016 219308
rect 244922 219328 244978 219337
rect 220266 219263 220322 219272
rect 248328 219302 248380 219308
rect 249432 219360 249484 219366
rect 249432 219302 249484 219308
rect 260748 219360 260800 219366
rect 260748 219302 260800 219308
rect 244922 219263 244978 219272
rect 9864 132932 9916 132938
rect 9864 132874 9916 132880
rect 20720 120760 20772 120766
rect 129004 120760 129056 120766
rect 43534 120728 43590 120737
rect 20720 120702 20772 120708
rect 10074 120006 10456 120034
rect 16698 120006 16804 120034
rect 10428 117978 10456 120006
rect 16776 118590 16804 120006
rect 16764 118584 16816 118590
rect 16764 118526 16816 118532
rect 10416 117972 10468 117978
rect 10416 117914 10468 117920
rect 15200 112396 15252 112402
rect 15200 112338 15252 112344
rect 9862 112024 9918 112033
rect 9862 111959 9918 111968
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 9876 3602 9904 111959
rect 15212 109956 15240 112338
rect 20732 109342 20760 120702
rect 43194 120686 43534 120714
rect 96434 120728 96490 120737
rect 96186 120686 96434 120714
rect 43534 120663 43590 120672
rect 103150 120728 103206 120737
rect 102810 120686 103150 120714
rect 96434 120663 96490 120672
rect 116398 120728 116454 120737
rect 116058 120686 116398 120714
rect 103150 120663 103206 120672
rect 216128 120760 216180 120766
rect 129056 120708 129306 120714
rect 129004 120702 129306 120708
rect 216128 120702 216180 120708
rect 129016 120686 129306 120702
rect 116398 120663 116454 120672
rect 29748 120142 29946 120170
rect 56244 120142 56442 120170
rect 155604 120142 155802 120170
rect 162228 120142 162426 120170
rect 195348 120142 195546 120170
rect 23032 120006 23322 120034
rect 23032 118658 23060 120006
rect 23020 118652 23072 118658
rect 23020 118594 23072 118600
rect 23032 117366 23060 118594
rect 29748 117881 29776 120142
rect 34978 120048 35034 120057
rect 38750 120048 38806 120057
rect 36570 120006 36676 120034
rect 34978 119983 35034 119992
rect 34992 119474 35020 119983
rect 35162 119912 35218 119921
rect 35162 119847 35218 119856
rect 35176 119474 35204 119847
rect 35346 119504 35402 119513
rect 34980 119468 35032 119474
rect 34980 119410 35032 119416
rect 35164 119468 35216 119474
rect 35346 119439 35348 119448
rect 35164 119410 35216 119416
rect 35400 119439 35402 119448
rect 35348 119410 35400 119416
rect 34886 119368 34942 119377
rect 34886 119303 34942 119312
rect 34900 119270 34928 119303
rect 34888 119264 34940 119270
rect 34888 119206 34940 119212
rect 34610 119096 34666 119105
rect 34610 119031 34612 119040
rect 34664 119031 34666 119040
rect 34612 119002 34664 119008
rect 34794 118960 34850 118969
rect 34794 118895 34850 118904
rect 34808 118862 34836 118895
rect 34796 118856 34848 118862
rect 34888 118856 34940 118862
rect 34796 118798 34848 118804
rect 34886 118824 34888 118833
rect 35164 118856 35216 118862
rect 34940 118824 34942 118833
rect 35164 118798 35216 118804
rect 34886 118759 34942 118768
rect 29734 117872 29790 117881
rect 29734 117807 29790 117816
rect 22100 117360 22152 117366
rect 22100 117302 22152 117308
rect 23020 117360 23072 117366
rect 23020 117302 23072 117308
rect 22112 109750 22140 117302
rect 32494 113928 32550 113937
rect 32494 113863 32496 113872
rect 32548 113863 32550 113872
rect 32496 113834 32548 113840
rect 28448 112600 28500 112606
rect 28448 112542 28500 112548
rect 28460 109956 28488 112542
rect 35070 112024 35126 112033
rect 35070 111959 35126 111968
rect 35084 109956 35112 111959
rect 35176 110702 35204 118798
rect 36648 117473 36676 120006
rect 49818 120006 49924 120034
rect 38750 119983 38806 119992
rect 38764 119474 38792 119983
rect 38752 119468 38804 119474
rect 38752 119410 38804 119416
rect 38844 119264 38896 119270
rect 38844 119206 38896 119212
rect 48134 119232 48190 119241
rect 38856 119105 38884 119206
rect 48134 119167 48190 119176
rect 38842 119096 38898 119105
rect 48148 119066 48176 119167
rect 38842 119031 38898 119040
rect 48136 119060 48188 119066
rect 48136 119002 48188 119008
rect 49896 118561 49924 120006
rect 56244 118658 56272 120142
rect 63498 120048 63554 120057
rect 62776 120006 63066 120034
rect 56232 118652 56284 118658
rect 56232 118594 56284 118600
rect 49882 118552 49938 118561
rect 49882 118487 49938 118496
rect 49896 117473 49924 118487
rect 56244 118153 56272 118594
rect 56230 118144 56286 118153
rect 56230 118079 56286 118088
rect 62776 117473 62804 120006
rect 63498 119983 63554 119992
rect 63682 120048 63738 120057
rect 69690 120006 70072 120034
rect 76314 120006 76420 120034
rect 82938 120006 83044 120034
rect 63682 119983 63738 119992
rect 63512 119542 63540 119983
rect 63500 119536 63552 119542
rect 63500 119478 63552 119484
rect 63696 119474 63724 119983
rect 63684 119468 63736 119474
rect 63684 119410 63736 119416
rect 64052 119468 64104 119474
rect 64052 119410 64104 119416
rect 64064 119377 64092 119410
rect 64050 119368 64106 119377
rect 64050 119303 64106 119312
rect 70044 117638 70072 120006
rect 76392 118153 76420 120006
rect 76378 118144 76434 118153
rect 76378 118079 76434 118088
rect 70032 117632 70084 117638
rect 70032 117574 70084 117580
rect 83016 117473 83044 120006
rect 89272 120006 89562 120034
rect 109144 120006 109434 120034
rect 122682 120006 122788 120034
rect 135930 120006 136036 120034
rect 36634 117464 36690 117473
rect 36634 117399 36690 117408
rect 49882 117464 49938 117473
rect 49882 117399 49938 117408
rect 62762 117464 62818 117473
rect 62762 117399 62818 117408
rect 83002 117464 83058 117473
rect 83002 117399 83058 117408
rect 89272 117366 89300 120006
rect 109144 118425 109172 120006
rect 109130 118416 109186 118425
rect 109130 118351 109186 118360
rect 122760 118114 122788 120006
rect 122196 118108 122248 118114
rect 122196 118050 122248 118056
rect 122748 118108 122800 118114
rect 122748 118050 122800 118056
rect 122208 117881 122236 118050
rect 122194 117872 122250 117881
rect 122194 117807 122250 117816
rect 136008 117473 136036 120006
rect 142356 120006 142554 120034
rect 149178 120006 149560 120034
rect 142356 118153 142384 120006
rect 145656 119468 145708 119474
rect 145656 119410 145708 119416
rect 145668 119105 145696 119410
rect 145748 119332 145800 119338
rect 145748 119274 145800 119280
rect 145654 119096 145710 119105
rect 145654 119031 145710 119040
rect 145668 118998 145696 119031
rect 145656 118992 145708 118998
rect 145656 118934 145708 118940
rect 145760 118833 145788 119274
rect 145746 118824 145802 118833
rect 145746 118759 145802 118768
rect 142342 118144 142398 118153
rect 142342 118079 142398 118088
rect 149532 117473 149560 120006
rect 155604 118590 155632 120142
rect 161018 120048 161074 120057
rect 161018 119983 161074 119992
rect 161032 119270 161060 119983
rect 161020 119264 161072 119270
rect 161020 119206 161072 119212
rect 157522 119096 157578 119105
rect 157522 119031 157578 119040
rect 157536 118998 157564 119031
rect 157524 118992 157576 118998
rect 157524 118934 157576 118940
rect 155592 118584 155644 118590
rect 155592 118526 155644 118532
rect 155604 117473 155632 118526
rect 162228 118522 162256 120142
rect 172702 120048 172758 120057
rect 168760 120006 169050 120034
rect 162490 119912 162546 119921
rect 162490 119847 162546 119856
rect 162504 119762 162532 119847
rect 162412 119734 162532 119762
rect 162412 119406 162440 119734
rect 162400 119400 162452 119406
rect 162400 119342 162452 119348
rect 162412 118862 162440 119342
rect 168104 118992 168156 118998
rect 168104 118934 168156 118940
rect 162400 118856 162452 118862
rect 162400 118798 162452 118804
rect 162216 118516 162268 118522
rect 162216 118458 162268 118464
rect 162228 117473 162256 118458
rect 135994 117464 136050 117473
rect 135994 117399 136050 117408
rect 149518 117464 149574 117473
rect 149518 117399 149574 117408
rect 155590 117464 155646 117473
rect 155590 117399 155646 117408
rect 162214 117464 162270 117473
rect 162214 117399 162270 117408
rect 89260 117360 89312 117366
rect 89260 117302 89312 117308
rect 106464 117360 106516 117366
rect 106464 117302 106516 117308
rect 69386 114472 69442 114481
rect 69386 114407 69442 114416
rect 69400 113422 69428 114407
rect 89272 114034 89300 117302
rect 89260 114028 89312 114034
rect 89260 113970 89312 113976
rect 69388 113416 69440 113422
rect 69388 113358 69440 113364
rect 81440 112532 81492 112538
rect 81440 112474 81492 112480
rect 48320 112464 48372 112470
rect 48320 112406 48372 112412
rect 41694 112024 41750 112033
rect 41694 111959 41750 111968
rect 35164 110696 35216 110702
rect 35164 110638 35216 110644
rect 41708 109956 41736 111959
rect 48332 109956 48360 112406
rect 61566 112160 61622 112169
rect 61566 112095 61622 112104
rect 68190 112160 68246 112169
rect 68190 112095 68246 112104
rect 54942 112024 54998 112033
rect 54942 111959 54998 111968
rect 54956 109956 54984 111959
rect 61580 109956 61608 112095
rect 68204 109956 68232 112095
rect 74814 112024 74870 112033
rect 74814 111959 74870 111968
rect 74828 109956 74856 111959
rect 81452 109956 81480 112474
rect 88062 112024 88118 112033
rect 88062 111959 88118 111968
rect 94686 112024 94742 112033
rect 94686 111959 94742 111968
rect 101310 112024 101366 112033
rect 101310 111959 101366 111968
rect 22100 109744 22152 109750
rect 22100 109686 22152 109692
rect 88076 109426 88104 111959
rect 94700 109956 94728 111959
rect 96896 110764 96948 110770
rect 96896 110706 96948 110712
rect 96908 110673 96936 110706
rect 96894 110664 96950 110673
rect 96894 110599 96950 110608
rect 101324 109956 101352 111959
rect 106476 111314 106504 117302
rect 160926 112840 160982 112849
rect 121184 112804 121236 112810
rect 160926 112775 160982 112784
rect 121184 112746 121236 112752
rect 107934 112568 107990 112577
rect 107934 112503 107990 112512
rect 106464 111308 106516 111314
rect 106464 111250 106516 111256
rect 106476 110770 106504 111250
rect 106464 110764 106516 110770
rect 106464 110706 106516 110712
rect 107948 109956 107976 112503
rect 115110 112160 115166 112169
rect 115110 112095 115166 112104
rect 115124 111926 115152 112095
rect 114560 111920 114612 111926
rect 114560 111862 114612 111868
rect 115112 111920 115164 111926
rect 115112 111862 115164 111868
rect 114572 109956 114600 111862
rect 121196 109956 121224 112746
rect 127808 112736 127860 112742
rect 127808 112678 127860 112684
rect 127820 109956 127848 112678
rect 141054 112568 141110 112577
rect 141054 112503 141110 112512
rect 134430 112160 134486 112169
rect 134430 112095 134486 112104
rect 132774 111616 132830 111625
rect 132774 111551 132776 111560
rect 132828 111551 132830 111560
rect 132776 111522 132828 111528
rect 134444 109956 134472 112095
rect 135720 111580 135772 111586
rect 135720 111522 135772 111528
rect 135732 110945 135760 111522
rect 135718 110936 135774 110945
rect 135718 110871 135774 110880
rect 137192 110560 137244 110566
rect 137190 110528 137192 110537
rect 137244 110528 137246 110537
rect 137190 110463 137246 110472
rect 141068 109956 141096 112503
rect 147678 112160 147734 112169
rect 147678 112095 147734 112104
rect 154302 112160 154358 112169
rect 154302 112095 154358 112104
rect 147692 109956 147720 112095
rect 154316 109956 154344 112095
rect 160940 109956 160968 112775
rect 162412 111314 162440 118798
rect 167550 112840 167606 112849
rect 167550 112775 167606 112784
rect 162400 111308 162452 111314
rect 162400 111250 162452 111256
rect 167564 109956 167592 112775
rect 168116 111654 168144 118934
rect 168760 118289 168788 120006
rect 175674 120006 175964 120034
rect 182298 120006 182680 120034
rect 188922 120006 189028 120034
rect 172702 119983 172758 119992
rect 172716 119270 172744 119983
rect 172704 119264 172756 119270
rect 172704 119206 172756 119212
rect 168746 118280 168802 118289
rect 168746 118215 168802 118224
rect 175936 117910 175964 120006
rect 179328 118924 179380 118930
rect 179328 118866 179380 118872
rect 175924 117904 175976 117910
rect 175924 117846 175976 117852
rect 175936 117473 175964 117846
rect 175922 117464 175978 117473
rect 175922 117399 175978 117408
rect 174174 111888 174230 111897
rect 174174 111823 174230 111832
rect 168104 111648 168156 111654
rect 168104 111590 168156 111596
rect 168116 110770 168144 111590
rect 168380 111308 168432 111314
rect 168380 111250 168432 111256
rect 168392 110809 168420 111250
rect 170218 111208 170274 111217
rect 170218 111143 170274 111152
rect 168378 110800 168434 110809
rect 168104 110764 168156 110770
rect 168378 110735 168380 110744
rect 168104 110706 168156 110712
rect 168432 110735 168434 110744
rect 168380 110706 168432 110712
rect 168104 110628 168156 110634
rect 168104 110570 168156 110576
rect 168116 110537 168144 110570
rect 170232 110566 170260 111143
rect 170220 110560 170272 110566
rect 168102 110528 168158 110537
rect 170220 110502 170272 110508
rect 168102 110463 168158 110472
rect 174188 109956 174216 111823
rect 179340 111353 179368 118866
rect 180892 118856 180944 118862
rect 180892 118798 180944 118804
rect 180798 112296 180854 112305
rect 180798 112231 180854 112240
rect 180614 111752 180670 111761
rect 180614 111687 180670 111696
rect 179510 111480 179566 111489
rect 179510 111415 179566 111424
rect 179326 111344 179382 111353
rect 179326 111279 179382 111288
rect 179340 111110 179368 111279
rect 179328 111104 179380 111110
rect 179328 111046 179380 111052
rect 179524 110566 179552 111415
rect 179880 111104 179932 111110
rect 179880 111046 179932 111052
rect 179892 110702 179920 111046
rect 180628 110770 180656 111687
rect 180616 110764 180668 110770
rect 180616 110706 180668 110712
rect 179880 110696 179932 110702
rect 179880 110638 179932 110644
rect 179512 110560 179564 110566
rect 179512 110502 179564 110508
rect 180812 109970 180840 112231
rect 180904 110702 180932 118798
rect 182652 117473 182680 120006
rect 189000 118289 189028 120006
rect 188986 118280 189042 118289
rect 188986 118215 189042 118224
rect 189000 117473 189028 118215
rect 195348 117842 195376 120142
rect 202170 120006 202276 120034
rect 208794 120006 209176 120034
rect 215418 120006 215524 120034
rect 202248 118386 202276 120006
rect 202236 118380 202288 118386
rect 202236 118322 202288 118328
rect 195336 117836 195388 117842
rect 195336 117778 195388 117784
rect 195348 117473 195376 117778
rect 202248 117473 202276 118322
rect 209148 118182 209176 120006
rect 215496 118318 215524 120006
rect 215758 119776 215814 119785
rect 215758 119711 215814 119720
rect 215574 119640 215630 119649
rect 215574 119575 215630 119584
rect 215588 119474 215616 119575
rect 215772 119474 215800 119711
rect 216034 119504 216090 119513
rect 215576 119468 215628 119474
rect 215576 119410 215628 119416
rect 215760 119468 215812 119474
rect 215760 119410 215812 119416
rect 215852 119468 215904 119474
rect 216140 119474 216168 120702
rect 248538 120698 248920 120714
rect 248538 120692 248932 120698
rect 248538 120686 248880 120692
rect 248880 120634 248932 120640
rect 299664 120692 299716 120698
rect 299664 120634 299716 120640
rect 221832 120148 221884 120154
rect 221832 120090 221884 120096
rect 216588 119672 216640 119678
rect 216588 119614 216640 119620
rect 216034 119439 216090 119448
rect 216128 119468 216180 119474
rect 215852 119410 215904 119416
rect 215864 119105 215892 119410
rect 216048 119406 216076 119439
rect 216128 119410 216180 119416
rect 216036 119400 216088 119406
rect 216036 119342 216088 119348
rect 216600 119105 216628 119614
rect 215850 119096 215906 119105
rect 215850 119031 215906 119040
rect 216586 119096 216642 119105
rect 216586 119031 216642 119040
rect 221844 118694 221872 120090
rect 222042 120006 222148 120034
rect 228666 120006 228864 120034
rect 235290 120006 235672 120034
rect 221844 118666 222056 118694
rect 215484 118312 215536 118318
rect 215484 118254 215536 118260
rect 209136 118176 209188 118182
rect 209134 118144 209136 118153
rect 209188 118144 209190 118153
rect 209134 118079 209190 118088
rect 182638 117464 182694 117473
rect 182638 117399 182694 117408
rect 188986 117464 189042 117473
rect 188986 117399 189042 117408
rect 195334 117464 195390 117473
rect 195334 117399 195390 117408
rect 202234 117464 202290 117473
rect 202234 117399 202290 117408
rect 209504 116612 209556 116618
rect 209504 116554 209556 116560
rect 209516 115802 209544 116554
rect 209870 115832 209926 115841
rect 209504 115796 209556 115802
rect 209870 115767 209926 115776
rect 209504 115738 209556 115744
rect 209884 115666 209912 115767
rect 209872 115660 209924 115666
rect 209872 115602 209924 115608
rect 209688 115592 209740 115598
rect 209688 115534 209740 115540
rect 187422 113112 187478 113121
rect 187422 113047 187478 113056
rect 194046 113112 194102 113121
rect 194046 113047 194102 113056
rect 183468 111716 183520 111722
rect 183468 111658 183520 111664
rect 181258 111616 181314 111625
rect 181258 111551 181314 111560
rect 181272 110702 181300 111551
rect 181352 111376 181404 111382
rect 183480 111353 183508 111658
rect 182638 111344 182694 111353
rect 181404 111324 181668 111330
rect 181352 111318 181668 111324
rect 181364 111314 181668 111318
rect 181364 111308 181680 111314
rect 181364 111302 181628 111308
rect 182638 111279 182694 111288
rect 183466 111344 183522 111353
rect 183466 111279 183522 111288
rect 181628 111250 181680 111256
rect 182088 111240 182140 111246
rect 181810 111208 181866 111217
rect 182088 111182 182140 111188
rect 181810 111143 181812 111152
rect 181864 111143 181866 111152
rect 181812 111114 181864 111120
rect 182100 110702 182128 111182
rect 182652 110770 182680 111279
rect 182824 111240 182876 111246
rect 183190 111208 183246 111217
rect 182876 111188 183140 111194
rect 182824 111182 183140 111188
rect 182836 111166 183140 111182
rect 183112 110974 183140 111166
rect 183190 111143 183246 111152
rect 183204 111042 183232 111143
rect 183192 111036 183244 111042
rect 183192 110978 183244 110984
rect 183100 110968 183152 110974
rect 183100 110910 183152 110916
rect 182640 110764 182692 110770
rect 182640 110706 182692 110712
rect 180892 110696 180944 110702
rect 180892 110638 180944 110644
rect 181260 110696 181312 110702
rect 181260 110638 181312 110644
rect 182088 110696 182140 110702
rect 182088 110638 182140 110644
rect 182652 110537 182680 110706
rect 182638 110528 182694 110537
rect 182638 110463 182694 110472
rect 180812 109956 180932 109970
rect 187436 109956 187464 113047
rect 190460 110560 190512 110566
rect 190458 110528 190460 110537
rect 190512 110528 190514 110537
rect 190458 110463 190514 110472
rect 194060 109956 194088 113047
rect 200670 112704 200726 112713
rect 200670 112639 200726 112648
rect 194508 111648 194560 111654
rect 194560 111596 194640 111602
rect 194508 111590 194640 111596
rect 194520 111574 194640 111590
rect 194414 111072 194470 111081
rect 194414 111007 194470 111016
rect 194428 110770 194456 111007
rect 194612 110770 194640 111574
rect 194324 110764 194376 110770
rect 194324 110706 194376 110712
rect 194416 110764 194468 110770
rect 194416 110706 194468 110712
rect 194600 110764 194652 110770
rect 194600 110706 194652 110712
rect 194692 110764 194744 110770
rect 194692 110706 194744 110712
rect 194336 110650 194364 110706
rect 194704 110650 194732 110706
rect 194336 110622 194732 110650
rect 200684 109956 200712 112639
rect 207294 111888 207350 111897
rect 207294 111823 207350 111832
rect 202524 110906 203104 110922
rect 202512 110900 203116 110906
rect 202564 110894 203064 110900
rect 202512 110842 202564 110848
rect 203064 110842 203116 110848
rect 207308 109956 207336 111823
rect 209700 111450 209728 115534
rect 220542 113112 220598 113121
rect 220542 113047 220598 113056
rect 213918 112704 213974 112713
rect 213918 112639 213974 112648
rect 213642 111480 213698 111489
rect 209688 111444 209740 111450
rect 213642 111415 213698 111424
rect 209688 111386 209740 111392
rect 213656 111246 213684 111415
rect 213644 111240 213696 111246
rect 213644 111182 213696 111188
rect 213932 109956 213960 112639
rect 220556 111994 220584 113047
rect 220544 111988 220596 111994
rect 220544 111930 220596 111936
rect 214564 111580 214616 111586
rect 214564 111522 214616 111528
rect 214470 111344 214526 111353
rect 214470 111279 214526 111288
rect 214484 110770 214512 111279
rect 214576 110945 214604 111522
rect 214654 111072 214710 111081
rect 214654 111007 214710 111016
rect 214562 110936 214618 110945
rect 214562 110871 214618 110880
rect 214668 110770 214696 111007
rect 214746 110936 214802 110945
rect 214746 110871 214802 110880
rect 214380 110764 214432 110770
rect 214380 110706 214432 110712
rect 214472 110764 214524 110770
rect 214472 110706 214524 110712
rect 214656 110764 214708 110770
rect 214656 110706 214708 110712
rect 214392 110650 214420 110706
rect 214392 110622 214512 110650
rect 214484 110566 214512 110622
rect 214380 110560 214432 110566
rect 214380 110502 214432 110508
rect 214472 110560 214524 110566
rect 214760 110514 214788 110871
rect 214472 110502 214524 110508
rect 214392 110378 214420 110502
rect 214576 110486 214788 110514
rect 214576 110378 214604 110486
rect 214392 110350 214604 110378
rect 220556 109956 220584 111930
rect 222028 111246 222056 118666
rect 222120 118318 222148 120006
rect 222108 118312 222160 118318
rect 222108 118254 222160 118260
rect 228836 118250 228864 120006
rect 235644 118561 235672 120006
rect 241716 120006 241914 120034
rect 239140 119610 239352 119626
rect 239128 119604 239364 119610
rect 239180 119598 239312 119604
rect 239128 119546 239180 119552
rect 239312 119546 239364 119552
rect 239404 119536 239456 119542
rect 239404 119478 239456 119484
rect 238760 119468 238812 119474
rect 238760 119410 238812 119416
rect 238852 119468 238904 119474
rect 238852 119410 238904 119416
rect 238772 119241 238800 119410
rect 238758 119232 238814 119241
rect 238758 119167 238814 119176
rect 238772 119066 238800 119167
rect 238760 119060 238812 119066
rect 238760 119002 238812 119008
rect 238864 118930 238892 119410
rect 239036 119400 239088 119406
rect 239312 119400 239364 119406
rect 239088 119348 239312 119354
rect 239036 119342 239364 119348
rect 239048 119326 239352 119342
rect 238944 119264 238996 119270
rect 239416 119218 239444 119478
rect 238996 119212 239444 119218
rect 238944 119206 239444 119212
rect 238956 119190 239444 119206
rect 238852 118924 238904 118930
rect 238852 118866 238904 118872
rect 235630 118552 235686 118561
rect 235630 118487 235686 118496
rect 228824 118244 228876 118250
rect 228824 118186 228876 118192
rect 228836 117473 228864 118186
rect 235644 117473 235672 118487
rect 241716 118289 241744 120006
rect 248512 119400 248564 119406
rect 248512 119342 248564 119348
rect 248236 119264 248288 119270
rect 248524 119218 248552 119342
rect 248288 119212 248552 119218
rect 248236 119206 248552 119212
rect 248248 119190 248552 119206
rect 241702 118280 241758 118289
rect 241702 118215 241758 118224
rect 241716 117473 241744 118215
rect 248892 118017 248920 120634
rect 254872 120006 255162 120034
rect 261496 120006 261786 120034
rect 268410 120006 268516 120034
rect 253940 119672 253992 119678
rect 253938 119640 253940 119649
rect 254492 119672 254544 119678
rect 253992 119640 253994 119649
rect 253938 119575 253994 119584
rect 254490 119640 254492 119649
rect 254544 119640 254546 119649
rect 254490 119575 254546 119584
rect 254216 119468 254268 119474
rect 254216 119410 254268 119416
rect 254228 119377 254256 119410
rect 254214 119368 254270 119377
rect 254214 119303 254270 119312
rect 254872 118425 254900 120006
rect 261496 118697 261524 120006
rect 261482 118688 261538 118697
rect 261482 118623 261538 118632
rect 254858 118416 254914 118425
rect 254858 118351 254914 118360
rect 268488 118153 268516 120006
rect 274652 120006 275034 120034
rect 281658 120006 282040 120034
rect 268474 118144 268530 118153
rect 268474 118079 268530 118088
rect 248878 118008 248934 118017
rect 248878 117943 248934 117952
rect 228822 117464 228878 117473
rect 228822 117399 228878 117408
rect 235630 117464 235686 117473
rect 235630 117399 235686 117408
rect 241702 117464 241758 117473
rect 241702 117399 241758 117408
rect 227166 113112 227222 113121
rect 227166 113047 227222 113056
rect 273258 113112 273314 113121
rect 273258 113047 273314 113056
rect 222384 111376 222436 111382
rect 222384 111318 222436 111324
rect 221924 111240 221976 111246
rect 221924 111182 221976 111188
rect 222016 111240 222068 111246
rect 222396 111217 222424 111318
rect 222016 111182 222068 111188
rect 222382 111208 222438 111217
rect 221936 110650 221964 111182
rect 222028 110770 222056 111182
rect 222382 111143 222438 111152
rect 222396 110770 222424 111143
rect 222016 110764 222068 110770
rect 222016 110706 222068 110712
rect 222200 110764 222252 110770
rect 222200 110706 222252 110712
rect 222384 110764 222436 110770
rect 222384 110706 222436 110712
rect 222568 110764 222620 110770
rect 222568 110706 222620 110712
rect 222108 110696 222160 110702
rect 221936 110644 222108 110650
rect 221936 110638 222160 110644
rect 221936 110622 222148 110638
rect 222212 110537 222240 110706
rect 222580 110650 222608 110706
rect 222396 110622 222608 110650
rect 222396 110566 222424 110622
rect 222384 110560 222436 110566
rect 222198 110528 222254 110537
rect 222384 110502 222436 110508
rect 222198 110463 222254 110472
rect 227180 109956 227208 113047
rect 273272 113014 273300 113047
rect 273260 113008 273312 113014
rect 273260 112950 273312 112956
rect 260288 112940 260340 112946
rect 260288 112882 260340 112888
rect 247038 112432 247094 112441
rect 247038 112367 247094 112376
rect 233790 112024 233846 112033
rect 233790 111959 233846 111968
rect 231858 111208 231914 111217
rect 231858 111143 231860 111152
rect 231912 111143 231914 111152
rect 231860 111114 231912 111120
rect 233804 109956 233832 111959
rect 240414 111888 240470 111897
rect 240414 111823 240470 111832
rect 240428 109956 240456 111823
rect 247052 109956 247080 112367
rect 253662 111888 253718 111897
rect 253662 111823 253718 111832
rect 253676 109956 253704 111823
rect 260300 109956 260328 112882
rect 266912 112872 266964 112878
rect 266912 112814 266964 112820
rect 266924 109956 266952 112814
rect 273166 110664 273222 110673
rect 273166 110599 273222 110608
rect 273180 110566 273208 110599
rect 273168 110560 273220 110566
rect 273168 110502 273220 110508
rect 273272 109970 273300 112950
rect 274180 111036 274232 111042
rect 274180 110978 274232 110984
rect 274192 110922 274220 110978
rect 273456 110906 274220 110922
rect 274652 110906 274680 120006
rect 282012 118454 282040 120006
rect 287992 120006 288282 120034
rect 294906 120006 295196 120034
rect 282000 118448 282052 118454
rect 282000 118390 282052 118396
rect 282012 117473 282040 118390
rect 281998 117464 282054 117473
rect 281998 117399 282054 117408
rect 287992 117337 288020 120006
rect 290462 119912 290518 119921
rect 290462 119847 290518 119856
rect 290476 119542 290504 119847
rect 290568 119610 290780 119626
rect 290556 119604 290792 119610
rect 290608 119598 290740 119604
rect 290556 119546 290608 119552
rect 290740 119546 290792 119552
rect 289912 119536 289964 119542
rect 289726 119504 289782 119513
rect 290464 119536 290516 119542
rect 289964 119484 290412 119490
rect 289912 119478 290412 119484
rect 290464 119478 290516 119484
rect 292118 119504 292174 119513
rect 289924 119462 290412 119478
rect 289726 119439 289728 119448
rect 289780 119439 289782 119448
rect 289728 119410 289780 119416
rect 290384 119406 290412 119462
rect 290372 119400 290424 119406
rect 290372 119342 290424 119348
rect 290476 119354 290504 119478
rect 292118 119439 292174 119448
rect 292132 119406 292160 119439
rect 292120 119400 292172 119406
rect 290476 119326 290780 119354
rect 292120 119342 292172 119348
rect 290752 119134 290780 119326
rect 290740 119128 290792 119134
rect 290740 119070 290792 119076
rect 295168 117774 295196 120006
rect 295156 117768 295208 117774
rect 295154 117736 295156 117745
rect 295208 117736 295210 117745
rect 295154 117671 295210 117680
rect 287978 117328 288034 117337
rect 287978 117263 288034 117272
rect 286782 112568 286838 112577
rect 286782 112503 286838 112512
rect 280158 111888 280214 111897
rect 280158 111823 280214 111832
rect 273444 110900 274220 110906
rect 273496 110894 274220 110900
rect 274640 110900 274692 110906
rect 273444 110842 273496 110848
rect 274640 110842 274692 110848
rect 273810 110800 273866 110809
rect 273810 110735 273866 110744
rect 273824 110702 273852 110735
rect 273444 110696 273496 110702
rect 273444 110638 273496 110644
rect 273628 110696 273680 110702
rect 273628 110638 273680 110644
rect 273812 110696 273864 110702
rect 273812 110638 273864 110644
rect 273456 110362 273484 110638
rect 273640 110537 273668 110638
rect 273626 110528 273682 110537
rect 273626 110463 273682 110472
rect 273444 110356 273496 110362
rect 273444 110298 273496 110304
rect 180826 109942 180932 109956
rect 273272 109942 273562 109970
rect 280172 109956 280200 111823
rect 286796 109956 286824 112503
rect 293408 112192 293460 112198
rect 293408 112134 293460 112140
rect 293420 111897 293448 112134
rect 293406 111888 293462 111897
rect 293406 111823 293462 111832
rect 293420 109956 293448 111823
rect 299676 109970 299704 120634
rect 301530 120006 301636 120034
rect 308154 120006 308536 120034
rect 301608 117706 301636 120006
rect 308312 119672 308364 119678
rect 307680 119620 308312 119626
rect 307680 119614 308364 119620
rect 307680 119610 308352 119614
rect 307668 119604 308352 119610
rect 307720 119598 308352 119604
rect 307668 119546 307720 119552
rect 308508 118046 308536 120006
rect 308496 118040 308548 118046
rect 308496 117982 308548 117988
rect 301596 117700 301648 117706
rect 301596 117642 301648 117648
rect 299676 109942 300058 109970
rect 88154 109440 88210 109449
rect 88076 109412 88154 109426
rect 88090 109398 88154 109412
rect 88154 109375 88210 109384
rect 180904 109342 180932 109942
rect 20720 109336 20772 109342
rect 20720 109278 20772 109284
rect 21548 109336 21600 109342
rect 180892 109336 180944 109342
rect 21600 109284 21850 109290
rect 21548 109278 21850 109284
rect 180892 109278 180944 109284
rect 21560 109262 21850 109278
rect 310072 67386 310100 255954
rect 310256 176186 310284 267854
rect 310428 256420 310480 256426
rect 310428 256362 310480 256368
rect 310440 256018 310468 256362
rect 310428 256012 310480 256018
rect 310428 255954 310480 255960
rect 310612 220040 310664 220046
rect 310612 219982 310664 219988
rect 310336 219768 310388 219774
rect 310336 219710 310388 219716
rect 310348 184006 310376 219710
rect 310520 217660 310572 217666
rect 310520 217602 310572 217608
rect 310532 210458 310560 217602
rect 310520 210452 310572 210458
rect 310520 210394 310572 210400
rect 310336 184000 310388 184006
rect 310336 183942 310388 183948
rect 310348 183666 310376 183942
rect 310336 183660 310388 183666
rect 310336 183602 310388 183608
rect 310624 183598 310652 219982
rect 310716 183666 310744 271118
rect 310808 224398 310836 334222
rect 311072 334212 311124 334218
rect 311072 334154 311124 334160
rect 311084 295662 311112 334154
rect 311072 295656 311124 295662
rect 311072 295598 311124 295604
rect 310796 224392 310848 224398
rect 310796 224334 310848 224340
rect 310980 219088 311032 219094
rect 310980 219030 311032 219036
rect 310796 218884 310848 218890
rect 310796 218826 310848 218832
rect 310808 183734 310836 218826
rect 310888 218748 310940 218754
rect 310888 218690 310940 218696
rect 310796 183728 310848 183734
rect 310796 183670 310848 183676
rect 310704 183660 310756 183666
rect 310704 183602 310756 183608
rect 310612 183592 310664 183598
rect 310612 183534 310664 183540
rect 310704 178560 310756 178566
rect 310704 178502 310756 178508
rect 310520 178288 310572 178294
rect 310520 178230 310572 178236
rect 310428 178220 310480 178226
rect 310428 178162 310480 178168
rect 310244 176180 310296 176186
rect 310244 176122 310296 176128
rect 310256 175642 310284 176122
rect 310244 175636 310296 175642
rect 310244 175578 310296 175584
rect 310256 113422 310284 175578
rect 310440 119610 310468 178162
rect 310428 119604 310480 119610
rect 310428 119546 310480 119552
rect 310428 117632 310480 117638
rect 310428 117574 310480 117580
rect 310244 113416 310296 113422
rect 310244 113358 310296 113364
rect 310336 111172 310388 111178
rect 310336 111114 310388 111120
rect 310060 67380 310112 67386
rect 310060 67322 310112 67328
rect 310348 45554 310376 111114
rect 310164 45526 310376 45554
rect 310164 44946 310192 45526
rect 310152 44940 310204 44946
rect 310152 44882 310204 44888
rect 310164 25362 310192 44882
rect 310440 44878 310468 117574
rect 310428 44872 310480 44878
rect 310428 44814 310480 44820
rect 310244 44736 310296 44742
rect 310244 44678 310296 44684
rect 310152 25356 310204 25362
rect 310152 25298 310204 25304
rect 29642 10704 29698 10713
rect 49882 10704 49938 10713
rect 29698 10676 29946 10690
rect 29698 10662 29960 10676
rect 49818 10662 49882 10690
rect 29642 10639 29698 10648
rect 10060 7546 10088 10132
rect 16684 8294 16712 10132
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 23308 8226 23336 10132
rect 23296 8220 23348 8226
rect 23296 8162 23348 8168
rect 23308 7614 23336 8162
rect 29932 7682 29960 10662
rect 49882 10639 49938 10648
rect 56138 10704 56194 10713
rect 62762 10704 62818 10713
rect 56194 10662 56442 10690
rect 56138 10639 56194 10648
rect 122378 10704 122434 10713
rect 62818 10676 63066 10690
rect 62818 10662 63080 10676
rect 62762 10639 62818 10648
rect 36556 9897 36584 10132
rect 36542 9888 36598 9897
rect 36542 9823 36598 9832
rect 35532 9376 35584 9382
rect 35530 9344 35532 9353
rect 35584 9344 35586 9353
rect 35530 9279 35586 9288
rect 36556 7750 36584 9823
rect 43180 8129 43208 10132
rect 43166 8120 43222 8129
rect 43166 8055 43222 8064
rect 42340 8016 42392 8022
rect 42340 7958 42392 7964
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 29920 7676 29972 7682
rect 29920 7618 29972 7624
rect 23296 7608 23348 7614
rect 23296 7550 23348 7556
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 21180 3664 21232 3670
rect 21180 3606 21232 3612
rect 39212 3664 39264 3670
rect 39212 3606 39264 3612
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 20 3392 72 3398
rect 20 3334 72 3340
rect 11978 3360 12034 3369
rect 32 480 60 3334
rect 11978 3295 12034 3304
rect 11992 480 12020 3295
rect 21192 480 21220 3606
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24136 480 24164 3538
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 36266 3496 36322 3505
rect 33336 480 33364 3470
rect 36266 3431 36322 3440
rect 36280 480 36308 3431
rect 39224 480 39252 3606
rect 42352 480 42380 7958
rect 63052 7818 63080 10662
rect 155498 10704 155554 10713
rect 122434 10662 122682 10690
rect 122378 10639 122434 10648
rect 162122 10704 162178 10713
rect 155554 10662 155802 10690
rect 155498 10639 155554 10648
rect 175922 10704 175978 10713
rect 162178 10662 162426 10690
rect 175674 10662 175922 10690
rect 162122 10639 162178 10648
rect 182638 10704 182694 10713
rect 182298 10676 182638 10690
rect 175922 10639 175978 10648
rect 182284 10662 182638 10676
rect 147956 10464 148008 10470
rect 147956 10406 148008 10412
rect 116768 10396 116820 10402
rect 116768 10338 116820 10344
rect 65154 9480 65210 9489
rect 65154 9415 65156 9424
rect 65208 9415 65210 9424
rect 66166 9480 66222 9489
rect 66166 9415 66222 9424
rect 65156 9386 65208 9392
rect 66180 9217 66208 9415
rect 66166 9208 66222 9217
rect 66166 9143 66222 9152
rect 63040 7812 63092 7818
rect 63040 7754 63092 7760
rect 69676 7478 69704 10132
rect 72240 9376 72292 9382
rect 72240 9318 72292 9324
rect 69664 7472 69716 7478
rect 69664 7414 69716 7420
rect 54484 5364 54536 5370
rect 54484 5306 54536 5312
rect 51354 3496 51410 3505
rect 51354 3431 51410 3440
rect 45284 3188 45336 3194
rect 45284 3130 45336 3136
rect 45296 480 45324 3130
rect 51368 480 51396 3431
rect 54496 480 54524 5306
rect 60556 5296 60608 5302
rect 60556 5238 60608 5244
rect 60568 480 60596 5238
rect 69572 3800 69624 3806
rect 69572 3742 69624 3748
rect 63500 3596 63552 3602
rect 63500 3538 63552 3544
rect 63512 480 63540 3538
rect 69584 480 69612 3742
rect 72252 3534 72280 9318
rect 76300 8265 76328 10132
rect 82924 9897 82952 10132
rect 82910 9888 82966 9897
rect 82910 9823 82966 9832
rect 77300 9648 77352 9654
rect 77298 9616 77300 9625
rect 78588 9648 78640 9654
rect 77352 9616 77354 9625
rect 77116 9580 77168 9586
rect 77298 9551 77354 9560
rect 77850 9616 77906 9625
rect 77850 9551 77852 9560
rect 77116 9522 77168 9528
rect 77904 9551 77906 9560
rect 78586 9616 78588 9625
rect 78640 9616 78642 9625
rect 78586 9551 78642 9560
rect 78864 9580 78916 9586
rect 77852 9522 77904 9528
rect 78864 9522 78916 9528
rect 79048 9580 79100 9586
rect 79048 9522 79100 9528
rect 77128 8945 77156 9522
rect 77944 9376 77996 9382
rect 77942 9344 77944 9353
rect 78876 9353 78904 9522
rect 79060 9489 79088 9522
rect 79232 9512 79284 9518
rect 79046 9480 79102 9489
rect 79046 9415 79102 9424
rect 79230 9480 79232 9489
rect 79284 9480 79286 9489
rect 79230 9415 79286 9424
rect 77996 9344 77998 9353
rect 77942 9279 77998 9288
rect 78862 9344 78918 9353
rect 78862 9279 78918 9288
rect 77114 8936 77170 8945
rect 77114 8871 77170 8880
rect 76286 8256 76342 8265
rect 76286 8191 76342 8200
rect 82924 7993 82952 9823
rect 88432 9580 88484 9586
rect 88432 9522 88484 9528
rect 88616 9580 88668 9586
rect 88616 9522 88668 9528
rect 88340 9444 88392 9450
rect 88340 9386 88392 9392
rect 88352 8537 88380 9386
rect 88444 8945 88472 9522
rect 88430 8936 88486 8945
rect 88430 8871 88486 8880
rect 88628 8809 88656 9522
rect 88614 8800 88670 8809
rect 88614 8735 88670 8744
rect 88338 8528 88394 8537
rect 88338 8463 88394 8472
rect 82910 7984 82966 7993
rect 82910 7919 82966 7928
rect 89548 7886 89576 10132
rect 95146 9616 95202 9625
rect 95146 9551 95148 9560
rect 95200 9551 95202 9560
rect 95148 9522 95200 9528
rect 96172 7993 96200 10132
rect 98828 9376 98880 9382
rect 98828 9318 98880 9324
rect 96158 7984 96214 7993
rect 96158 7919 96214 7928
rect 88524 7880 88576 7886
rect 88524 7822 88576 7828
rect 89536 7880 89588 7886
rect 89536 7822 89588 7828
rect 78588 7676 78640 7682
rect 78588 7618 78640 7624
rect 75644 7608 75696 7614
rect 75644 7550 75696 7556
rect 72240 3528 72292 3534
rect 72240 3470 72292 3476
rect 72698 3496 72754 3505
rect 72698 3431 72754 3440
rect 72712 480 72740 3431
rect 75656 480 75684 7550
rect 78600 480 78628 7618
rect 88536 4826 88564 7822
rect 88524 4820 88576 4826
rect 88524 4762 88576 4768
rect 98840 4078 98868 9318
rect 102796 7857 102824 10132
rect 109420 8129 109448 10132
rect 109406 8120 109462 8129
rect 109406 8055 109462 8064
rect 116044 7993 116072 10132
rect 116490 9616 116546 9625
rect 116780 9586 116808 10338
rect 116490 9551 116492 9560
rect 116544 9551 116546 9560
rect 116584 9580 116636 9586
rect 116492 9522 116544 9528
rect 116584 9522 116636 9528
rect 116768 9580 116820 9586
rect 116768 9522 116820 9528
rect 116596 8974 116624 9522
rect 116584 8968 116636 8974
rect 116584 8910 116636 8916
rect 117044 8968 117096 8974
rect 117044 8910 117096 8916
rect 116030 7984 116086 7993
rect 116030 7919 116086 7928
rect 102782 7848 102838 7857
rect 102782 7783 102838 7792
rect 98828 4072 98880 4078
rect 98828 4014 98880 4020
rect 102874 4040 102930 4049
rect 102874 3975 102930 3984
rect 100114 3768 100170 3777
rect 100114 3703 100170 3712
rect 100128 3505 100156 3703
rect 99930 3496 99986 3505
rect 99930 3431 99986 3440
rect 100114 3496 100170 3505
rect 100114 3431 100170 3440
rect 99944 480 99972 3431
rect 102888 480 102916 3975
rect 106002 3768 106058 3777
rect 106002 3703 106058 3712
rect 108948 3732 109000 3738
rect 106016 480 106044 3703
rect 108948 3674 109000 3680
rect 108960 480 108988 3674
rect 117056 3398 117084 8910
rect 129292 8158 129320 10132
rect 135916 9897 135944 10132
rect 142264 10118 142554 10146
rect 142264 9897 142292 10118
rect 135902 9888 135958 9897
rect 135902 9823 135958 9832
rect 142250 9888 142306 9897
rect 142250 9823 142306 9832
rect 129280 8152 129332 8158
rect 129280 8094 129332 8100
rect 135916 7954 135944 9823
rect 147968 9586 147996 10406
rect 151268 10328 151320 10334
rect 151268 10270 151320 10276
rect 149518 10160 149574 10169
rect 149178 10132 149518 10146
rect 149164 10118 149518 10132
rect 147956 9580 148008 9586
rect 147956 9522 148008 9528
rect 148048 9580 148100 9586
rect 148048 9522 148100 9528
rect 147772 9376 147824 9382
rect 147772 9318 147824 9324
rect 147784 9042 147812 9318
rect 148060 9081 148088 9522
rect 148046 9072 148102 9081
rect 147772 9036 147824 9042
rect 148046 9007 148102 9016
rect 147772 8978 147824 8984
rect 149164 8090 149192 10118
rect 149518 10095 149574 10104
rect 151280 9722 151308 10270
rect 168656 9920 168708 9926
rect 168656 9862 168708 9868
rect 168470 9752 168526 9761
rect 151268 9716 151320 9722
rect 168668 9722 168696 9862
rect 168930 9752 168986 9761
rect 168470 9687 168526 9696
rect 168656 9716 168708 9722
rect 151268 9658 151320 9664
rect 150992 9580 151044 9586
rect 150992 9522 151044 9528
rect 152556 9580 152608 9586
rect 152556 9522 152608 9528
rect 151004 8906 151032 9522
rect 152568 8945 152596 9522
rect 152554 8936 152610 8945
rect 150992 8900 151044 8906
rect 152554 8871 152610 8880
rect 150992 8842 151044 8848
rect 168484 8566 168512 9687
rect 168930 9687 168932 9696
rect 168656 9658 168708 9664
rect 168984 9687 168986 9696
rect 168932 9658 168984 9664
rect 168840 9648 168892 9654
rect 168746 9616 168802 9625
rect 168892 9596 168972 9602
rect 168840 9590 168972 9596
rect 168852 9586 168972 9590
rect 168852 9580 168984 9586
rect 168852 9574 168932 9580
rect 168746 9551 168748 9560
rect 168800 9551 168802 9560
rect 168748 9522 168800 9528
rect 168932 9522 168984 9528
rect 168656 9512 168708 9518
rect 168656 9454 168708 9460
rect 168668 8566 168696 9454
rect 168472 8560 168524 8566
rect 168472 8502 168524 8508
rect 168656 8560 168708 8566
rect 168656 8502 168708 8508
rect 149152 8084 149204 8090
rect 149152 8026 149204 8032
rect 135904 7948 135956 7954
rect 135904 7890 135956 7896
rect 168668 7886 168696 8502
rect 169036 8129 169064 10132
rect 169116 9920 169168 9926
rect 169116 9862 169168 9868
rect 169128 9692 169156 9862
rect 169116 9686 169168 9692
rect 169116 9628 169168 9634
rect 169298 9616 169354 9625
rect 169298 9551 169300 9560
rect 169352 9551 169354 9560
rect 169300 9522 169352 9528
rect 170140 9302 170444 9330
rect 170140 9178 170168 9302
rect 170312 9240 170364 9246
rect 170232 9188 170312 9194
rect 170232 9182 170364 9188
rect 170128 9172 170180 9178
rect 170128 9114 170180 9120
rect 170232 9166 170352 9182
rect 170416 9178 170444 9302
rect 170404 9172 170456 9178
rect 170232 9110 170260 9166
rect 170404 9114 170456 9120
rect 170220 9104 170272 9110
rect 170220 9046 170272 9052
rect 169022 8120 169078 8129
rect 169022 8055 169078 8064
rect 168656 7880 168708 7886
rect 168656 7822 168708 7828
rect 182284 6914 182312 10662
rect 188986 10704 189042 10713
rect 188922 10662 188986 10690
rect 182638 10639 182694 10648
rect 188986 10639 189042 10648
rect 195242 10704 195298 10713
rect 202234 10704 202290 10713
rect 195298 10662 195546 10690
rect 202170 10662 202234 10690
rect 195242 10639 195298 10648
rect 208858 10704 208914 10713
rect 208794 10662 208858 10690
rect 202234 10639 202290 10648
rect 208858 10639 208914 10648
rect 228362 10704 228418 10713
rect 235630 10704 235686 10713
rect 228418 10662 228666 10690
rect 235290 10662 235630 10690
rect 228362 10639 228418 10648
rect 248878 10704 248934 10713
rect 248538 10676 248878 10690
rect 235630 10639 235686 10648
rect 248524 10662 248878 10676
rect 239956 10600 240008 10606
rect 239956 10542 240008 10548
rect 185766 9616 185822 9625
rect 185766 9551 185822 9560
rect 185780 9382 185808 9551
rect 185768 9376 185820 9382
rect 185768 9318 185820 9324
rect 215404 8022 215432 10132
rect 222028 8158 222056 10132
rect 239968 9722 239996 10542
rect 244648 10532 244700 10538
rect 244648 10474 244700 10480
rect 244554 10296 244610 10305
rect 244554 10231 244610 10240
rect 241702 10160 241758 10169
rect 241758 10132 241914 10146
rect 241758 10118 241928 10132
rect 241702 10095 241758 10104
rect 239956 9716 240008 9722
rect 239956 9658 240008 9664
rect 239864 9580 239916 9586
rect 239864 9522 239916 9528
rect 240048 9580 240100 9586
rect 240048 9522 240100 9528
rect 239876 9081 239904 9522
rect 240060 9217 240088 9522
rect 240046 9208 240102 9217
rect 240046 9143 240102 9152
rect 239862 9072 239918 9081
rect 239862 9007 239918 9016
rect 239876 8673 239904 9007
rect 239862 8664 239918 8673
rect 239862 8599 239918 8608
rect 240060 8498 240088 9143
rect 240048 8492 240100 8498
rect 240048 8434 240100 8440
rect 222016 8152 222068 8158
rect 222016 8094 222068 8100
rect 215392 8016 215444 8022
rect 215392 7958 215444 7964
rect 241900 7614 241928 10118
rect 244568 9586 244596 10231
rect 244660 9586 244688 10474
rect 248144 9716 248196 9722
rect 248144 9658 248196 9664
rect 244556 9580 244608 9586
rect 244556 9522 244608 9528
rect 244648 9580 244700 9586
rect 244648 9522 244700 9528
rect 244280 9512 244332 9518
rect 244280 9454 244332 9460
rect 244292 8809 244320 9454
rect 244278 8800 244334 8809
rect 244278 8735 244334 8744
rect 244660 8430 244688 9522
rect 248156 9489 248184 9658
rect 248142 9480 248198 9489
rect 248142 9415 248198 9424
rect 244648 8424 244700 8430
rect 244648 8366 244700 8372
rect 241888 7608 241940 7614
rect 241888 7550 241940 7556
rect 248524 6914 248552 10662
rect 248878 10639 248934 10648
rect 254858 10704 254914 10713
rect 261482 10704 261538 10713
rect 254914 10662 255162 10690
rect 254858 10639 254914 10648
rect 268750 10704 268806 10713
rect 261538 10662 261786 10690
rect 261852 10668 261904 10674
rect 261482 10639 261538 10648
rect 268410 10662 268750 10690
rect 268750 10639 268806 10648
rect 274730 10704 274786 10713
rect 281998 10704 282054 10713
rect 274786 10662 275034 10690
rect 281658 10662 281998 10690
rect 274730 10639 274786 10648
rect 281998 10639 282054 10648
rect 287978 10704 288034 10713
rect 294602 10704 294658 10713
rect 288034 10662 288282 10690
rect 287978 10639 288034 10648
rect 294658 10662 294906 10690
rect 294602 10639 294658 10648
rect 261852 10610 261904 10616
rect 261760 9512 261812 9518
rect 261312 9460 261760 9466
rect 261312 9454 261812 9460
rect 261312 9438 261800 9454
rect 261312 9382 261340 9438
rect 261300 9376 261352 9382
rect 261300 9318 261352 9324
rect 261484 9376 261536 9382
rect 261864 9330 261892 10610
rect 310164 10606 310192 25298
rect 310152 10600 310204 10606
rect 310152 10542 310204 10548
rect 272340 9716 272392 9722
rect 272340 9658 272392 9664
rect 277768 9716 277820 9722
rect 277768 9658 277820 9664
rect 272156 9648 272208 9654
rect 272062 9616 272118 9625
rect 270684 9580 270736 9586
rect 270684 9522 270736 9528
rect 270868 9580 270920 9586
rect 272156 9590 272208 9596
rect 272062 9551 272118 9560
rect 270868 9522 270920 9528
rect 261536 9324 261892 9330
rect 261484 9318 261892 9324
rect 261496 9302 261892 9318
rect 270696 9217 270724 9522
rect 270880 9353 270908 9522
rect 272076 9518 272104 9551
rect 270960 9512 271012 9518
rect 270960 9454 271012 9460
rect 272064 9512 272116 9518
rect 272064 9454 272116 9460
rect 270866 9344 270922 9353
rect 270866 9279 270922 9288
rect 270682 9208 270738 9217
rect 270682 9143 270738 9152
rect 270972 8945 271000 9454
rect 271328 9444 271380 9450
rect 271328 9386 271380 9392
rect 270958 8936 271014 8945
rect 270958 8871 271014 8880
rect 271340 8430 271368 9386
rect 272168 9081 272196 9590
rect 272154 9072 272210 9081
rect 272154 9007 272210 9016
rect 271328 8424 271380 8430
rect 272352 8401 272380 9658
rect 277780 9625 277808 9658
rect 278136 9648 278188 9654
rect 273166 9616 273222 9625
rect 277766 9616 277822 9625
rect 273166 9551 273168 9560
rect 273220 9551 273222 9560
rect 277676 9580 277728 9586
rect 273168 9522 273220 9528
rect 278136 9590 278188 9596
rect 277766 9551 277822 9560
rect 277676 9522 277728 9528
rect 273442 9480 273498 9489
rect 277688 9466 277716 9522
rect 273442 9415 273498 9424
rect 277504 9438 277716 9466
rect 273456 9382 273484 9415
rect 277504 9382 277532 9438
rect 273444 9376 273496 9382
rect 277492 9376 277544 9382
rect 273444 9318 273496 9324
rect 273810 9344 273866 9353
rect 277492 9318 277544 9324
rect 277584 9376 277636 9382
rect 277584 9318 277636 9324
rect 273810 9279 273866 9288
rect 273824 8634 273852 9279
rect 277596 8945 277624 9318
rect 278044 9240 278096 9246
rect 277688 9188 278044 9194
rect 277688 9182 278096 9188
rect 277688 9166 278084 9182
rect 277582 8936 277638 8945
rect 277582 8871 277638 8880
rect 277688 8634 277716 9166
rect 278148 9081 278176 9590
rect 280896 9308 280948 9314
rect 280896 9250 280948 9256
rect 280908 9110 280936 9250
rect 280896 9104 280948 9110
rect 278134 9072 278190 9081
rect 280896 9046 280948 9052
rect 282092 9104 282144 9110
rect 282092 9046 282144 9052
rect 278134 9007 278190 9016
rect 282104 8650 282132 9046
rect 273812 8628 273864 8634
rect 273812 8570 273864 8576
rect 277676 8628 277728 8634
rect 282104 8622 282316 8650
rect 277676 8570 277728 8576
rect 282288 8566 282316 8622
rect 282276 8560 282328 8566
rect 282276 8502 282328 8508
rect 271328 8366 271380 8372
rect 272338 8392 272394 8401
rect 272338 8327 272394 8336
rect 301516 8294 301544 10132
rect 301504 8288 301556 8294
rect 301504 8230 301556 8236
rect 308140 8226 308168 10132
rect 308128 8220 308180 8226
rect 308128 8162 308180 8168
rect 278596 7812 278648 7818
rect 278596 7754 278648 7760
rect 272524 7744 272576 7750
rect 272524 7686 272576 7692
rect 182192 6886 182312 6914
rect 248432 6886 248552 6914
rect 148324 4820 148376 4826
rect 148324 4762 148376 4768
rect 124034 3768 124090 3777
rect 124034 3703 124090 3712
rect 117044 3392 117096 3398
rect 117044 3334 117096 3340
rect 124048 480 124076 3703
rect 145380 3392 145432 3398
rect 145380 3334 145432 3340
rect 142250 3088 142306 3097
rect 142250 3023 142306 3032
rect 142264 480 142292 3023
rect 145392 480 145420 3334
rect 148336 480 148364 4762
rect 178682 4040 178738 4049
rect 178682 3975 178738 3984
rect 151450 3904 151506 3913
rect 151450 3839 151506 3848
rect 151464 480 151492 3839
rect 175554 3632 175610 3641
rect 175554 3567 175610 3576
rect 157340 3324 157392 3330
rect 157340 3266 157392 3272
rect 157352 480 157380 3266
rect 172612 3256 172664 3262
rect 169482 3224 169538 3233
rect 172612 3198 172664 3204
rect 169482 3159 169538 3168
rect 169496 480 169524 3159
rect 172624 480 172652 3198
rect 175568 480 175596 3567
rect 178696 480 178724 3975
rect 182192 3194 182220 6886
rect 205916 5092 205968 5098
rect 205916 5034 205968 5040
rect 193772 4004 193824 4010
rect 193772 3946 193824 3952
rect 182180 3188 182232 3194
rect 182180 3130 182232 3136
rect 193784 3126 193812 3946
rect 193772 3120 193824 3126
rect 193772 3062 193824 3068
rect 193784 480 193812 3062
rect 205928 480 205956 5034
rect 208860 4004 208912 4010
rect 208860 3946 208912 3952
rect 208872 480 208900 3946
rect 233148 3936 233200 3942
rect 233148 3878 233200 3884
rect 211986 3768 212042 3777
rect 211986 3703 212042 3712
rect 212000 480 212028 3703
rect 221002 3496 221058 3505
rect 221002 3431 221058 3440
rect 214932 3188 214984 3194
rect 214932 3130 214984 3136
rect 214944 480 214972 3130
rect 221016 480 221044 3431
rect 230204 3052 230256 3058
rect 230204 2994 230256 3000
rect 230216 480 230244 2994
rect 233160 480 233188 3878
rect 236092 3868 236144 3874
rect 236092 3810 236144 3816
rect 236104 480 236132 3810
rect 242162 3632 242218 3641
rect 242162 3567 242218 3576
rect 242176 480 242204 3567
rect 248432 3126 248460 6886
rect 263506 4040 263562 4049
rect 263506 3975 263562 3984
rect 257436 3868 257488 3874
rect 257436 3810 257488 3816
rect 251362 3496 251418 3505
rect 251362 3431 251418 3440
rect 248420 3120 248472 3126
rect 248420 3062 248472 3068
rect 251376 480 251404 3431
rect 254308 2984 254360 2990
rect 254308 2926 254360 2932
rect 254320 480 254348 2926
rect 257448 480 257476 3810
rect 260380 2916 260432 2922
rect 260380 2858 260432 2864
rect 260392 480 260420 2858
rect 263520 480 263548 3975
rect 266450 3768 266506 3777
rect 266450 3703 266506 3712
rect 266464 480 266492 3703
rect 272536 480 272564 7686
rect 278608 480 278636 7754
rect 310256 7478 310284 44678
rect 310244 7472 310296 7478
rect 310244 7414 310296 7420
rect 293684 4072 293736 4078
rect 293684 4014 293736 4020
rect 302884 4072 302936 4078
rect 302884 4014 302936 4020
rect 281538 3632 281594 3641
rect 281538 3567 281594 3576
rect 281552 480 281580 3567
rect 287612 3120 287664 3126
rect 287612 3062 287664 3068
rect 284668 2848 284720 2854
rect 284668 2790 284720 2796
rect 284680 480 284708 2790
rect 287624 480 287652 3062
rect 293696 480 293724 4014
rect 302896 480 302924 4014
rect 310532 2990 310560 178230
rect 310716 178158 310744 178502
rect 310900 178362 310928 218690
rect 310888 178356 310940 178362
rect 310888 178298 310940 178304
rect 310704 178152 310756 178158
rect 310704 178094 310756 178100
rect 310716 176202 310744 178094
rect 310796 178084 310848 178090
rect 310796 178026 310848 178032
rect 310624 176174 310744 176202
rect 310624 120766 310652 176174
rect 310704 176044 310756 176050
rect 310704 175986 310756 175992
rect 310612 120760 310664 120766
rect 310612 120702 310664 120708
rect 310610 45928 310666 45937
rect 310610 45863 310666 45872
rect 310624 25362 310652 45863
rect 310612 25356 310664 25362
rect 310612 25298 310664 25304
rect 310716 9586 310744 175986
rect 310808 116618 310836 178026
rect 310992 176050 311020 219030
rect 311072 202156 311124 202162
rect 311072 202098 311124 202104
rect 310980 176044 311032 176050
rect 310980 175986 311032 175992
rect 311084 120834 311112 202098
rect 311072 120828 311124 120834
rect 311072 120770 311124 120776
rect 311176 119882 311204 549238
rect 311348 441652 311400 441658
rect 311348 441594 311400 441600
rect 311256 331424 311308 331430
rect 311256 331366 311308 331372
rect 311164 119876 311216 119882
rect 311164 119818 311216 119824
rect 310980 117700 311032 117706
rect 310980 117642 311032 117648
rect 310796 116612 310848 116618
rect 310796 116554 310848 116560
rect 310888 110628 310940 110634
rect 310888 110570 310940 110576
rect 310704 9580 310756 9586
rect 310704 9522 310756 9528
rect 310900 4078 310928 110570
rect 310992 8294 311020 117642
rect 311164 110560 311216 110566
rect 311164 110502 311216 110508
rect 310980 8288 311032 8294
rect 310980 8230 311032 8236
rect 310888 4072 310940 4078
rect 310888 4014 310940 4020
rect 311176 3058 311204 110502
rect 311268 3398 311296 331366
rect 311360 119746 311388 441594
rect 311820 426766 311848 616762
rect 313384 586226 313412 616762
rect 313568 615738 313596 619520
rect 315396 616684 315448 616690
rect 315396 616626 315448 616632
rect 314108 616412 314160 616418
rect 314108 616354 314160 616360
rect 314016 616004 314068 616010
rect 314016 615946 314068 615952
rect 313556 615732 313608 615738
rect 313556 615674 313608 615680
rect 313372 586220 313424 586226
rect 313372 586162 313424 586168
rect 313924 555144 313976 555150
rect 313924 555086 313976 555092
rect 311900 465248 311952 465254
rect 311900 465190 311952 465196
rect 311808 426760 311860 426766
rect 311808 426702 311860 426708
rect 311624 368960 311676 368966
rect 311624 368902 311676 368908
rect 311440 244384 311492 244390
rect 311440 244326 311492 244332
rect 311348 119740 311400 119746
rect 311348 119682 311400 119688
rect 311348 30728 311400 30734
rect 311348 30670 311400 30676
rect 311256 3392 311308 3398
rect 311256 3334 311308 3340
rect 311360 3194 311388 30670
rect 311452 3194 311480 244326
rect 311532 219020 311584 219026
rect 311532 218962 311584 218968
rect 311544 178294 311572 218962
rect 311636 183802 311664 368902
rect 311714 220144 311770 220153
rect 311714 220079 311770 220088
rect 311624 183796 311676 183802
rect 311624 183738 311676 183744
rect 311532 178288 311584 178294
rect 311532 178230 311584 178236
rect 311532 125996 311584 126002
rect 311532 125938 311584 125944
rect 311544 25294 311572 125938
rect 311624 118788 311676 118794
rect 311624 118730 311676 118736
rect 311636 36582 311664 118730
rect 311728 48278 311756 220079
rect 311808 218952 311860 218958
rect 311808 218894 311860 218900
rect 311820 202026 311848 218894
rect 311808 202020 311860 202026
rect 311808 201962 311860 201968
rect 311808 183660 311860 183666
rect 311808 183602 311860 183608
rect 311820 121786 311848 183602
rect 311808 121780 311860 121786
rect 311808 121722 311860 121728
rect 311716 48272 311768 48278
rect 311716 48214 311768 48220
rect 311912 45082 311940 465190
rect 312084 424516 312136 424522
rect 312084 424458 312136 424464
rect 312096 423706 312124 424458
rect 312084 423700 312136 423706
rect 312084 423642 312136 423648
rect 311992 383784 312044 383790
rect 311992 383726 312044 383732
rect 312004 120902 312032 383726
rect 312096 205193 312124 423642
rect 312176 401668 312228 401674
rect 312176 401610 312228 401616
rect 312082 205184 312138 205193
rect 312082 205119 312138 205128
rect 312188 185609 312216 401610
rect 312544 359168 312596 359174
rect 312544 359110 312596 359116
rect 312268 337748 312320 337754
rect 312268 337690 312320 337696
rect 312174 185600 312230 185609
rect 312174 185535 312230 185544
rect 312082 166016 312138 166025
rect 312082 165951 312138 165960
rect 311992 120896 312044 120902
rect 311992 120838 312044 120844
rect 311992 85536 312044 85542
rect 311990 85504 311992 85513
rect 312044 85504 312046 85513
rect 311990 85439 312046 85448
rect 311900 45076 311952 45082
rect 311900 45018 311952 45024
rect 311624 36576 311676 36582
rect 311624 36518 311676 36524
rect 311532 25288 311584 25294
rect 311532 25230 311584 25236
rect 311898 17912 311954 17921
rect 311898 17847 311954 17856
rect 311912 16969 311940 17847
rect 311898 16960 311954 16969
rect 311898 16895 311954 16904
rect 311912 6914 311940 16895
rect 312004 16574 312032 85439
rect 312096 56001 312124 165951
rect 312174 156224 312230 156233
rect 312174 156159 312230 156168
rect 312188 126002 312216 156159
rect 312280 146441 312308 337690
rect 312360 337544 312412 337550
rect 312360 337486 312412 337492
rect 312372 175817 312400 337486
rect 312452 289876 312504 289882
rect 312452 289818 312504 289824
rect 312464 214985 312492 289818
rect 312556 216850 312584 359110
rect 313832 319456 313884 319462
rect 313832 319398 313884 319404
rect 313188 219836 313240 219842
rect 313188 219778 313240 219784
rect 312544 216844 312596 216850
rect 312544 216786 312596 216792
rect 313200 216782 313228 219778
rect 313188 216776 313240 216782
rect 313188 216718 313240 216724
rect 312450 214976 312506 214985
rect 312450 214911 312506 214920
rect 312634 214976 312690 214985
rect 312634 214911 312690 214920
rect 312542 205184 312598 205193
rect 312542 205119 312598 205128
rect 312450 185600 312506 185609
rect 312450 185535 312506 185544
rect 312358 175808 312414 175817
rect 312358 175743 312414 175752
rect 312266 146432 312322 146441
rect 312266 146367 312322 146376
rect 312266 126848 312322 126857
rect 312266 126783 312322 126792
rect 312280 126342 312308 126783
rect 312268 126336 312320 126342
rect 312268 126278 312320 126284
rect 312176 125996 312228 126002
rect 312176 125938 312228 125944
rect 312082 55992 312138 56001
rect 312082 55927 312138 55936
rect 312280 17921 312308 126278
rect 312372 66201 312400 175743
rect 312464 75857 312492 185535
rect 312556 95169 312584 205119
rect 312648 105641 312676 214911
rect 313844 201482 313872 319398
rect 313832 201476 313884 201482
rect 313832 201418 313884 201424
rect 312910 195392 312966 195401
rect 312910 195327 312966 195336
rect 312726 146432 312782 146441
rect 312726 146367 312782 146376
rect 312740 107710 312768 146367
rect 312818 136640 312874 136649
rect 312818 136575 312874 136584
rect 312728 107704 312780 107710
rect 312728 107646 312780 107652
rect 312634 105632 312690 105641
rect 312634 105567 312690 105576
rect 312542 95160 312598 95169
rect 312542 95095 312598 95104
rect 312544 85808 312596 85814
rect 312544 85750 312596 85756
rect 312450 75848 312506 75857
rect 312450 75783 312506 75792
rect 312358 66192 312414 66201
rect 312358 66127 312414 66136
rect 312450 55992 312506 56001
rect 312450 55927 312506 55936
rect 312464 55894 312492 55927
rect 312452 55888 312504 55894
rect 312452 55830 312504 55836
rect 312556 27305 312584 85750
rect 312740 36718 312768 107646
rect 312832 85746 312860 136575
rect 312820 85740 312872 85746
rect 312820 85682 312872 85688
rect 312924 85542 312952 195327
rect 313832 142180 313884 142186
rect 313832 142122 313884 142128
rect 313740 119128 313792 119134
rect 313740 119070 313792 119076
rect 312912 85536 312964 85542
rect 312912 85478 312964 85484
rect 313752 57458 313780 119070
rect 313740 57452 313792 57458
rect 313740 57394 313792 57400
rect 312728 36712 312780 36718
rect 312726 36680 312728 36689
rect 312780 36680 312782 36689
rect 312636 36644 312688 36650
rect 312726 36615 312782 36624
rect 312636 36586 312688 36592
rect 312542 27296 312598 27305
rect 312542 27231 312598 27240
rect 312266 17912 312322 17921
rect 312266 17847 312322 17856
rect 312004 16546 312124 16574
rect 311912 6886 312032 6914
rect 311900 3392 311952 3398
rect 311900 3334 311952 3340
rect 311348 3188 311400 3194
rect 311348 3130 311400 3136
rect 311440 3188 311492 3194
rect 311440 3130 311492 3136
rect 311164 3052 311216 3058
rect 311164 2994 311216 3000
rect 310520 2984 310572 2990
rect 310520 2926 310572 2932
rect 311912 480 311940 3334
rect 312004 3330 312032 6886
rect 311992 3324 312044 3330
rect 311992 3266 312044 3272
rect 312096 2854 312124 16546
rect 312648 2922 312676 36586
rect 313844 3806 313872 142122
rect 313832 3800 313884 3806
rect 313832 3742 313884 3748
rect 313936 3505 313964 555086
rect 314028 63782 314056 615946
rect 314120 117094 314148 616354
rect 314200 599004 314252 599010
rect 314200 598946 314252 598952
rect 314212 119678 314240 598946
rect 314292 454368 314344 454374
rect 314292 454310 314344 454316
rect 314200 119672 314252 119678
rect 314200 119614 314252 119620
rect 314108 117088 314160 117094
rect 314108 117030 314160 117036
rect 314108 111036 314160 111042
rect 314108 110978 314160 110984
rect 314120 66638 314148 110978
rect 314108 66632 314160 66638
rect 314108 66574 314160 66580
rect 314016 63776 314068 63782
rect 314016 63718 314068 63724
rect 313922 3496 313978 3505
rect 313922 3431 313978 3440
rect 314304 2922 314332 454310
rect 315304 453280 315356 453286
rect 315304 453222 315356 453228
rect 314384 399968 314436 399974
rect 314384 399910 314436 399916
rect 314396 3330 314424 399910
rect 314568 365764 314620 365770
rect 314568 365706 314620 365712
rect 314476 321632 314528 321638
rect 314476 321574 314528 321580
rect 314488 46374 314516 321574
rect 314580 116686 314608 365706
rect 315120 248736 315172 248742
rect 315120 248678 315172 248684
rect 314568 116680 314620 116686
rect 314568 116622 314620 116628
rect 314476 46368 314528 46374
rect 314476 46310 314528 46316
rect 315132 3806 315160 248678
rect 315212 147552 315264 147558
rect 315212 147494 315264 147500
rect 315224 108594 315252 147494
rect 315212 108588 315264 108594
rect 315212 108530 315264 108536
rect 315316 4078 315344 453222
rect 315408 114918 315436 616626
rect 315764 469260 315816 469266
rect 315764 469202 315816 469208
rect 315488 267776 315540 267782
rect 315488 267718 315540 267724
rect 315396 114912 315448 114918
rect 315396 114854 315448 114860
rect 315396 110968 315448 110974
rect 315396 110910 315448 110916
rect 315408 59634 315436 110910
rect 315396 59628 315448 59634
rect 315396 59570 315448 59576
rect 315500 10674 315528 267718
rect 315776 240922 315804 469202
rect 316052 362574 316080 619534
rect 316512 619426 316540 619534
rect 316654 619520 316766 620960
rect 318812 619534 319484 619562
rect 316696 619426 316724 619520
rect 316512 619398 316724 619426
rect 316684 556708 316736 556714
rect 316684 556650 316736 556656
rect 316040 362568 316092 362574
rect 316040 362510 316092 362516
rect 315764 240916 315816 240922
rect 315764 240858 315816 240864
rect 315580 228064 315632 228070
rect 315580 228006 315632 228012
rect 315488 10668 315540 10674
rect 315488 10610 315540 10616
rect 315304 4072 315356 4078
rect 315304 4014 315356 4020
rect 315120 3800 315172 3806
rect 315120 3742 315172 3748
rect 314384 3324 314436 3330
rect 314384 3266 314436 3272
rect 314844 3052 314896 3058
rect 314844 2994 314896 3000
rect 312636 2916 312688 2922
rect 312636 2858 312688 2864
rect 314292 2916 314344 2922
rect 314292 2858 314344 2864
rect 312084 2848 312136 2854
rect 312084 2790 312136 2796
rect 314856 480 314884 2994
rect 315592 2990 315620 228006
rect 315672 220176 315724 220182
rect 315672 220118 315724 220124
rect 315684 15434 315712 220118
rect 315764 195016 315816 195022
rect 315764 194958 315816 194964
rect 315672 15428 315724 15434
rect 315672 15370 315724 15376
rect 315580 2984 315632 2990
rect 315580 2926 315632 2932
rect 315776 2854 315804 194958
rect 315948 161492 316000 161498
rect 315948 161434 316000 161440
rect 315960 3058 315988 161434
rect 316592 142860 316644 142866
rect 316592 142802 316644 142808
rect 316604 111110 316632 142802
rect 316696 112334 316724 556650
rect 316776 554804 316828 554810
rect 316776 554746 316828 554752
rect 316788 118114 316816 554746
rect 317328 510944 317380 510950
rect 317328 510886 317380 510892
rect 316868 407176 316920 407182
rect 316868 407118 316920 407124
rect 316776 118108 316828 118114
rect 316776 118050 316828 118056
rect 316880 117910 316908 407118
rect 316960 397588 317012 397594
rect 316960 397530 317012 397536
rect 316868 117904 316920 117910
rect 316868 117846 316920 117852
rect 316972 117842 317000 397530
rect 317052 383716 317104 383722
rect 317052 383658 317104 383664
rect 316960 117836 317012 117842
rect 316960 117778 317012 117784
rect 316684 112328 316736 112334
rect 316684 112270 316736 112276
rect 316592 111104 316644 111110
rect 316592 111046 316644 111052
rect 317064 107846 317092 383658
rect 317236 220244 317288 220250
rect 317236 220186 317288 220192
rect 317144 219700 317196 219706
rect 317144 219642 317196 219648
rect 317052 107840 317104 107846
rect 317052 107782 317104 107788
rect 317156 15910 317184 219642
rect 317248 107982 317276 220186
rect 317236 107976 317288 107982
rect 317236 107918 317288 107924
rect 317144 15904 317196 15910
rect 317144 15846 317196 15852
rect 317340 9586 317368 510886
rect 318064 414316 318116 414322
rect 318064 414258 318116 414264
rect 317696 260160 317748 260166
rect 317696 260102 317748 260108
rect 317708 118726 317736 260102
rect 317972 118992 318024 118998
rect 317972 118934 318024 118940
rect 317696 118720 317748 118726
rect 317696 118662 317748 118668
rect 317984 105126 318012 118934
rect 317972 105120 318024 105126
rect 317972 105062 318024 105068
rect 318076 84794 318104 414258
rect 318812 337550 318840 619534
rect 319456 619426 319484 619534
rect 319598 619520 319710 620960
rect 322726 619520 322838 620960
rect 325670 619520 325782 620960
rect 328614 619520 328726 620960
rect 331742 619520 331854 620960
rect 334686 619520 334798 620960
rect 337814 619520 337926 620960
rect 340758 619520 340870 620960
rect 343886 619520 343998 620960
rect 346830 619520 346942 620960
rect 349958 619520 350070 620960
rect 351932 619534 352788 619562
rect 319640 619426 319668 619520
rect 319456 619398 319668 619426
rect 322204 616616 322256 616622
rect 322204 616558 322256 616564
rect 319904 514888 319956 514894
rect 319904 514830 319956 514836
rect 319812 514820 319864 514826
rect 319812 514762 319864 514768
rect 318800 337544 318852 337550
rect 318800 337486 318852 337492
rect 318156 334076 318208 334082
rect 318156 334018 318208 334024
rect 318168 123078 318196 334018
rect 319824 260982 319852 514762
rect 319812 260976 319864 260982
rect 319812 260918 319864 260924
rect 319916 260914 319944 514830
rect 321468 282600 321520 282606
rect 321468 282542 321520 282548
rect 319904 260908 319956 260914
rect 319904 260850 319956 260856
rect 318524 220516 318576 220522
rect 318524 220458 318576 220464
rect 318246 220280 318302 220289
rect 318246 220215 318302 220224
rect 318156 123072 318208 123078
rect 318156 123014 318208 123020
rect 318156 119060 318208 119066
rect 318156 119002 318208 119008
rect 318064 84788 318116 84794
rect 318064 84730 318116 84736
rect 318168 57254 318196 119002
rect 318156 57248 318208 57254
rect 318156 57190 318208 57196
rect 318064 45824 318116 45830
rect 318064 45766 318116 45772
rect 317328 9580 317380 9586
rect 317328 9522 317380 9528
rect 318076 5234 318104 45766
rect 318260 15502 318288 220215
rect 318340 219972 318392 219978
rect 318340 219914 318392 219920
rect 318352 30326 318380 219914
rect 318432 219564 318484 219570
rect 318432 219506 318484 219512
rect 318340 30320 318392 30326
rect 318340 30262 318392 30268
rect 318444 30258 318472 219506
rect 318536 46102 318564 220458
rect 318708 220176 318760 220182
rect 318708 220118 318760 220124
rect 318720 219910 318748 220118
rect 318708 219904 318760 219910
rect 318708 219846 318760 219852
rect 318616 118856 318668 118862
rect 318616 118798 318668 118804
rect 318628 89894 318656 118798
rect 318616 89888 318668 89894
rect 318616 89830 318668 89836
rect 318524 46096 318576 46102
rect 318524 46038 318576 46044
rect 318720 46034 318748 219846
rect 321480 152658 321508 282542
rect 321928 257440 321980 257446
rect 321928 257382 321980 257388
rect 321468 152652 321520 152658
rect 321468 152594 321520 152600
rect 321376 151904 321428 151910
rect 321376 151846 321428 151852
rect 319444 130416 319496 130422
rect 319444 130358 319496 130364
rect 319456 112606 319484 130358
rect 319444 112600 319496 112606
rect 319444 112542 319496 112548
rect 320180 55888 320232 55894
rect 320180 55830 320232 55836
rect 318708 46028 318760 46034
rect 318708 45970 318760 45976
rect 318432 30252 318484 30258
rect 318432 30194 318484 30200
rect 318248 15496 318300 15502
rect 318248 15438 318300 15444
rect 320192 6914 320220 55830
rect 321388 31482 321416 151846
rect 321376 31476 321428 31482
rect 321376 31418 321428 31424
rect 320456 30320 320508 30326
rect 320456 30262 320508 30268
rect 320468 8702 320496 30262
rect 321480 8838 321508 152594
rect 321940 152046 321968 257382
rect 322216 200870 322244 616558
rect 328656 605834 328684 619520
rect 331784 616418 331812 619520
rect 331772 616412 331824 616418
rect 331772 616354 331824 616360
rect 334728 615602 334756 619520
rect 334716 615596 334768 615602
rect 334716 615538 334768 615544
rect 334728 615494 334756 615538
rect 328472 605806 328684 605834
rect 334636 615466 334756 615494
rect 337856 615494 337884 619520
rect 337856 615466 338068 615494
rect 325608 599072 325660 599078
rect 325608 599014 325660 599020
rect 325620 566030 325648 599014
rect 325608 566024 325660 566030
rect 325608 565966 325660 565972
rect 325792 566024 325844 566030
rect 325792 565966 325844 565972
rect 325516 565956 325568 565962
rect 325516 565898 325568 565904
rect 324964 507816 325016 507822
rect 324964 507758 325016 507764
rect 324976 507686 325004 507758
rect 324964 507680 325016 507686
rect 324964 507622 325016 507628
rect 324976 492046 325004 507622
rect 324964 492040 325016 492046
rect 324964 491982 325016 491988
rect 322296 383240 322348 383246
rect 322296 383182 322348 383188
rect 322204 200864 322256 200870
rect 322204 200806 322256 200812
rect 321928 152040 321980 152046
rect 321928 151982 321980 151988
rect 321652 151972 321704 151978
rect 321652 151914 321704 151920
rect 321664 121854 321692 151914
rect 321652 121848 321704 121854
rect 321652 121790 321704 121796
rect 321468 8832 321520 8838
rect 321468 8774 321520 8780
rect 320456 8696 320508 8702
rect 320456 8638 320508 8644
rect 320192 6886 320496 6914
rect 318064 5228 318116 5234
rect 318064 5170 318116 5176
rect 315948 3052 316000 3058
rect 315948 2994 316000 3000
rect 317972 3052 318024 3058
rect 317972 2994 318024 3000
rect 315764 2848 315816 2854
rect 315764 2790 315816 2796
rect 317984 480 318012 2994
rect 320468 490 320496 6886
rect 322308 3262 322336 383182
rect 325528 369102 325556 565898
rect 325804 410922 325832 565966
rect 327264 556980 327316 556986
rect 327264 556922 327316 556928
rect 326344 539300 326396 539306
rect 326344 539242 326396 539248
rect 326356 508026 326384 539242
rect 326344 508020 326396 508026
rect 326344 507962 326396 507968
rect 325792 410916 325844 410922
rect 325792 410858 325844 410864
rect 326528 397792 326580 397798
rect 326528 397734 326580 397740
rect 325516 369096 325568 369102
rect 325516 369038 325568 369044
rect 323584 353388 323636 353394
rect 323584 353330 323636 353336
rect 323596 152658 323624 353330
rect 324964 294024 325016 294030
rect 324964 293966 325016 293972
rect 324976 175234 325004 293966
rect 324964 175228 325016 175234
rect 324964 175170 325016 175176
rect 323584 152652 323636 152658
rect 323584 152594 323636 152600
rect 326540 5370 326568 397734
rect 326988 355360 327040 355366
rect 326988 355302 327040 355308
rect 326528 5364 326580 5370
rect 326528 5306 326580 5312
rect 322296 3256 322348 3262
rect 322296 3198 322348 3204
rect 320744 598 320956 626
rect 320744 490 320772 598
rect -10 -960 102 480
rect 2934 -960 3046 480
rect 5878 -960 5990 480
rect 9006 -960 9118 480
rect 11950 -960 12062 480
rect 15078 -960 15190 480
rect 18022 -960 18134 480
rect 21150 -960 21262 480
rect 24094 -960 24206 480
rect 27222 -960 27334 480
rect 30166 -960 30278 480
rect 33294 -960 33406 480
rect 36238 -960 36350 480
rect 39182 -960 39294 480
rect 42310 -960 42422 480
rect 45254 -960 45366 480
rect 48382 -960 48494 480
rect 51326 -960 51438 480
rect 54454 -960 54566 480
rect 57398 -960 57510 480
rect 60526 -960 60638 480
rect 63470 -960 63582 480
rect 66598 -960 66710 480
rect 69542 -960 69654 480
rect 72670 -960 72782 480
rect 75614 -960 75726 480
rect 78558 -960 78670 480
rect 81686 -960 81798 480
rect 84630 -960 84742 480
rect 87758 -960 87870 480
rect 90702 -960 90814 480
rect 93830 -960 93942 480
rect 96774 -960 96886 480
rect 99902 -960 100014 480
rect 102846 -960 102958 480
rect 105974 -960 106086 480
rect 108918 -960 109030 480
rect 112046 -960 112158 480
rect 114990 -960 115102 480
rect 117934 -960 118046 480
rect 121062 -960 121174 480
rect 124006 -960 124118 480
rect 127134 -960 127246 480
rect 130078 -960 130190 480
rect 133206 -960 133318 480
rect 136150 -960 136262 480
rect 139278 -960 139390 480
rect 142222 -960 142334 480
rect 145350 -960 145462 480
rect 148294 -960 148406 480
rect 151422 -960 151534 480
rect 154366 -960 154478 480
rect 157310 -960 157422 480
rect 160438 -960 160550 480
rect 163382 -960 163494 480
rect 166510 -960 166622 480
rect 169454 -960 169566 480
rect 172582 -960 172694 480
rect 175526 -960 175638 480
rect 178654 -960 178766 480
rect 181598 -960 181710 480
rect 184726 -960 184838 480
rect 187670 -960 187782 480
rect 190798 -960 190910 480
rect 193742 -960 193854 480
rect 196686 -960 196798 480
rect 199814 -960 199926 480
rect 202758 -960 202870 480
rect 205886 -960 205998 480
rect 208830 -960 208942 480
rect 211958 -960 212070 480
rect 214902 -960 215014 480
rect 218030 -960 218142 480
rect 220974 -960 221086 480
rect 224102 -960 224214 480
rect 227046 -960 227158 480
rect 230174 -960 230286 480
rect 233118 -960 233230 480
rect 236062 -960 236174 480
rect 239190 -960 239302 480
rect 242134 -960 242246 480
rect 245262 -960 245374 480
rect 248206 -960 248318 480
rect 251334 -960 251446 480
rect 254278 -960 254390 480
rect 257406 -960 257518 480
rect 260350 -960 260462 480
rect 263478 -960 263590 480
rect 266422 -960 266534 480
rect 269550 -960 269662 480
rect 272494 -960 272606 480
rect 275438 -960 275550 480
rect 278566 -960 278678 480
rect 281510 -960 281622 480
rect 284638 -960 284750 480
rect 287582 -960 287694 480
rect 290710 -960 290822 480
rect 293654 -960 293766 480
rect 296782 -960 296894 480
rect 299726 -960 299838 480
rect 302854 -960 302966 480
rect 305798 -960 305910 480
rect 308926 -960 309038 480
rect 311870 -960 311982 480
rect 314814 -960 314926 480
rect 317942 -960 318054 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 327000 480 327028 355302
rect 327276 111858 327304 556922
rect 328472 514010 328500 605806
rect 331220 599276 331272 599282
rect 331220 599218 331272 599224
rect 330852 554056 330904 554062
rect 330852 553998 330904 554004
rect 330864 542366 330892 553998
rect 330852 542360 330904 542366
rect 330852 542302 330904 542308
rect 328460 514004 328512 514010
rect 328460 513946 328512 513952
rect 327724 480616 327776 480622
rect 327724 480558 327776 480564
rect 327356 112328 327408 112334
rect 327356 112270 327408 112276
rect 327368 111858 327396 112270
rect 327264 111852 327316 111858
rect 327264 111794 327316 111800
rect 327356 111852 327408 111858
rect 327356 111794 327408 111800
rect 327736 85610 327764 480558
rect 328472 223038 328500 513946
rect 331232 423502 331260 599218
rect 331496 556844 331548 556850
rect 331496 556786 331548 556792
rect 331508 534682 331536 556786
rect 331496 534676 331548 534682
rect 331496 534618 331548 534624
rect 331312 534472 331364 534478
rect 331312 534414 331364 534420
rect 331220 423496 331272 423502
rect 331220 423438 331272 423444
rect 330484 392352 330536 392358
rect 330484 392294 330536 392300
rect 329748 280492 329800 280498
rect 329748 280434 329800 280440
rect 329760 227730 329788 280434
rect 329748 227724 329800 227730
rect 329748 227666 329800 227672
rect 328460 223032 328512 223038
rect 328460 222974 328512 222980
rect 328552 115592 328604 115598
rect 328552 115534 328604 115540
rect 328564 112266 328592 115534
rect 328552 112260 328604 112266
rect 328552 112202 328604 112208
rect 328276 112192 328328 112198
rect 328276 112134 328328 112140
rect 327908 112056 327960 112062
rect 327908 111998 327960 112004
rect 327920 103514 327948 111998
rect 327828 103486 327948 103514
rect 327724 85604 327776 85610
rect 327724 85546 327776 85552
rect 327828 78606 327856 103486
rect 327816 78600 327868 78606
rect 327816 78542 327868 78548
rect 328288 8430 328316 112134
rect 328564 111858 328592 112202
rect 328552 111852 328604 111858
rect 328552 111794 328604 111800
rect 328276 8424 328328 8430
rect 328276 8366 328328 8372
rect 330496 3262 330524 392294
rect 331232 260166 331260 423438
rect 331220 260160 331272 260166
rect 331220 260102 331272 260108
rect 331324 209774 331352 534414
rect 331508 534342 331536 534618
rect 331496 534336 331548 534342
rect 331496 534278 331548 534284
rect 331588 497888 331640 497894
rect 331588 497830 331640 497836
rect 331404 423564 331456 423570
rect 331404 423506 331456 423512
rect 331416 263974 331444 423506
rect 331496 423496 331548 423502
rect 331496 423438 331548 423444
rect 331508 410582 331536 423438
rect 331496 410576 331548 410582
rect 331496 410518 331548 410524
rect 331600 325106 331628 497830
rect 331680 478916 331732 478922
rect 331680 478858 331732 478864
rect 331692 423502 331720 478858
rect 334636 467498 334664 615466
rect 334900 607980 334952 607986
rect 334900 607922 334952 607928
rect 334716 607776 334768 607782
rect 334716 607718 334768 607724
rect 334728 543862 334756 607718
rect 334716 543856 334768 543862
rect 334716 543798 334768 543804
rect 334912 534478 334940 607922
rect 334900 534472 334952 534478
rect 334900 534414 334952 534420
rect 334624 467492 334676 467498
rect 334624 467434 334676 467440
rect 338040 463758 338068 615466
rect 343928 605834 343956 619520
rect 346492 615936 346544 615942
rect 346492 615878 346544 615884
rect 343652 605806 343956 605834
rect 343652 548554 343680 605806
rect 343640 548548 343692 548554
rect 343640 548490 343692 548496
rect 342444 531616 342496 531622
rect 342444 531558 342496 531564
rect 340880 466880 340932 466886
rect 340880 466822 340932 466828
rect 338028 463752 338080 463758
rect 338028 463694 338080 463700
rect 333520 451376 333572 451382
rect 333520 451318 333572 451324
rect 333532 446758 333560 451318
rect 333520 446752 333572 446758
rect 333520 446694 333572 446700
rect 331680 423496 331732 423502
rect 331680 423438 331732 423444
rect 331772 334212 331824 334218
rect 331772 334154 331824 334160
rect 331784 325106 331812 334154
rect 331588 325100 331640 325106
rect 331588 325042 331640 325048
rect 331772 325100 331824 325106
rect 331772 325042 331824 325048
rect 331404 263968 331456 263974
rect 331404 263910 331456 263916
rect 331232 209746 331352 209774
rect 331232 202842 331260 209746
rect 331220 202836 331272 202842
rect 331220 202778 331272 202784
rect 331232 201958 331260 202778
rect 331220 201952 331272 201958
rect 331220 201894 331272 201900
rect 331864 123616 331916 123622
rect 331864 123558 331916 123564
rect 331876 3398 331904 123558
rect 333060 7948 333112 7954
rect 333060 7890 333112 7896
rect 331864 3392 331916 3398
rect 331864 3334 331916 3340
rect 330484 3256 330536 3262
rect 330484 3198 330536 3204
rect 333072 480 333100 7890
rect 333532 3058 333560 446694
rect 336556 439816 336608 439822
rect 336556 439758 336608 439764
rect 334072 417580 334124 417586
rect 334072 417522 334124 417528
rect 334084 383858 334112 417522
rect 334348 417512 334400 417518
rect 334348 417454 334400 417460
rect 334072 383852 334124 383858
rect 334072 383794 334124 383800
rect 334084 373994 334112 383794
rect 333992 373966 334112 373994
rect 333992 267734 334020 373966
rect 333992 267706 334112 267734
rect 333980 256488 334032 256494
rect 333980 256430 334032 256436
rect 333992 256086 334020 256430
rect 333980 256080 334032 256086
rect 333980 256022 334032 256028
rect 334084 256018 334112 267706
rect 334360 256494 334388 417454
rect 335544 410644 335596 410650
rect 335544 410586 335596 410592
rect 334348 256488 334400 256494
rect 334348 256430 334400 256436
rect 334072 256012 334124 256018
rect 334072 255954 334124 255960
rect 335556 15366 335584 410586
rect 335636 369164 335688 369170
rect 335636 369106 335688 369112
rect 335648 15366 335676 369106
rect 336188 360256 336240 360262
rect 336188 360198 336240 360204
rect 336096 252000 336148 252006
rect 336096 251942 336148 251948
rect 335912 225004 335964 225010
rect 335912 224946 335964 224952
rect 335924 175982 335952 224946
rect 336108 176118 336136 251942
rect 336200 176186 336228 360198
rect 336568 176186 336596 439758
rect 338764 433356 338816 433362
rect 338764 433298 338816 433304
rect 338212 421252 338264 421258
rect 338212 421194 338264 421200
rect 337752 282192 337804 282198
rect 337752 282134 337804 282140
rect 336188 176180 336240 176186
rect 336188 176122 336240 176128
rect 336556 176180 336608 176186
rect 336556 176122 336608 176128
rect 336096 176112 336148 176118
rect 336096 176054 336148 176060
rect 335912 175976 335964 175982
rect 335912 175918 335964 175924
rect 337476 175840 337528 175846
rect 337476 175782 337528 175788
rect 337488 111858 337516 175782
rect 337476 111852 337528 111858
rect 337476 111794 337528 111800
rect 337764 78674 337792 282134
rect 338224 78674 338252 421194
rect 337752 78668 337804 78674
rect 337752 78610 337804 78616
rect 338212 78668 338264 78674
rect 338212 78610 338264 78616
rect 338028 78600 338080 78606
rect 338028 78542 338080 78548
rect 335544 15360 335596 15366
rect 335544 15302 335596 15308
rect 335636 15360 335688 15366
rect 335636 15302 335688 15308
rect 338040 3670 338068 78542
rect 338776 39846 338804 433298
rect 340892 291378 340920 466822
rect 342260 375624 342312 375630
rect 342260 375566 342312 375572
rect 342272 319122 342300 375566
rect 342260 319116 342312 319122
rect 342260 319058 342312 319064
rect 340972 318912 341024 318918
rect 340972 318854 341024 318860
rect 342076 318912 342128 318918
rect 342076 318854 342128 318860
rect 340880 291372 340932 291378
rect 340880 291314 340932 291320
rect 339960 260296 340012 260302
rect 339960 260238 340012 260244
rect 339316 78600 339368 78606
rect 339316 78542 339368 78548
rect 339328 67250 339356 78542
rect 339316 67244 339368 67250
rect 339316 67186 339368 67192
rect 339972 45966 340000 260238
rect 340420 220108 340472 220114
rect 340420 220050 340472 220056
rect 340432 216714 340460 220050
rect 340420 216708 340472 216714
rect 340420 216650 340472 216656
rect 339960 45960 340012 45966
rect 339960 45902 340012 45908
rect 338764 39840 338816 39846
rect 338764 39782 338816 39788
rect 339972 5030 340000 45902
rect 340420 45824 340472 45830
rect 340420 45766 340472 45772
rect 340432 8090 340460 45766
rect 340892 8498 340920 291314
rect 340984 119202 341012 318854
rect 341432 291372 341484 291378
rect 341432 291314 341484 291320
rect 341340 291304 341392 291310
rect 341340 291246 341392 291252
rect 341248 291236 341300 291242
rect 341248 291178 341300 291184
rect 341156 236224 341208 236230
rect 341156 236166 341208 236172
rect 340972 119196 341024 119202
rect 340972 119138 341024 119144
rect 341168 8974 341196 236166
rect 341260 220794 341288 291178
rect 341248 220788 341300 220794
rect 341248 220730 341300 220736
rect 341352 220454 341380 291246
rect 341340 220448 341392 220454
rect 341340 220390 341392 220396
rect 341444 111654 341472 291314
rect 342088 119746 342116 318854
rect 342352 236224 342404 236230
rect 342352 236166 342404 236172
rect 342076 119740 342128 119746
rect 342076 119682 342128 119688
rect 341432 111648 341484 111654
rect 341432 111590 341484 111596
rect 342364 10402 342392 236166
rect 342352 10396 342404 10402
rect 342352 10338 342404 10344
rect 341156 8968 341208 8974
rect 341156 8910 341208 8916
rect 340880 8492 340932 8498
rect 340880 8434 340932 8440
rect 340420 8084 340472 8090
rect 340420 8026 340472 8032
rect 342456 5302 342484 531558
rect 344284 470892 344336 470898
rect 344284 470834 344336 470840
rect 342904 409420 342956 409426
rect 342904 409362 342956 409368
rect 342536 319116 342588 319122
rect 342536 319058 342588 319064
rect 342548 236366 342576 319058
rect 342536 236360 342588 236366
rect 342536 236302 342588 236308
rect 342548 220590 342576 236302
rect 342536 220584 342588 220590
rect 342536 220526 342588 220532
rect 342916 59430 342944 409362
rect 344296 59498 344324 470834
rect 346504 387598 346532 615878
rect 351460 525224 351512 525230
rect 351460 525166 351512 525172
rect 351736 525224 351788 525230
rect 351736 525166 351788 525172
rect 349804 505164 349856 505170
rect 349804 505106 349856 505112
rect 346860 415472 346912 415478
rect 346860 415414 346912 415420
rect 346584 415404 346636 415410
rect 346584 415346 346636 415352
rect 346596 387598 346624 415346
rect 346872 387666 346900 415414
rect 346768 387660 346820 387666
rect 346768 387602 346820 387608
rect 346860 387660 346912 387666
rect 346860 387602 346912 387608
rect 346492 387592 346544 387598
rect 346492 387534 346544 387540
rect 346584 387592 346636 387598
rect 346584 387534 346636 387540
rect 346308 387456 346360 387462
rect 346308 387398 346360 387404
rect 344744 339244 344796 339250
rect 344744 339186 344796 339192
rect 344756 301510 344784 339186
rect 344928 339040 344980 339046
rect 344928 338982 344980 338988
rect 344744 301504 344796 301510
rect 344744 301446 344796 301452
rect 344756 301170 344784 301446
rect 344744 301164 344796 301170
rect 344744 301106 344796 301112
rect 344652 102196 344704 102202
rect 344652 102138 344704 102144
rect 344284 59492 344336 59498
rect 344284 59434 344336 59440
rect 342904 59424 342956 59430
rect 342904 59366 342956 59372
rect 343916 36168 343968 36174
rect 343916 36110 343968 36116
rect 343928 8566 343956 36110
rect 344664 12442 344692 102138
rect 344940 61266 344968 338982
rect 344928 61260 344980 61266
rect 344928 61202 344980 61208
rect 346320 36106 346348 387398
rect 346504 36378 346532 387534
rect 346780 113286 346808 387602
rect 346872 178566 346900 387602
rect 348424 322720 348476 322726
rect 348424 322662 348476 322668
rect 347044 258120 347096 258126
rect 347044 258062 347096 258068
rect 347056 225690 347084 258062
rect 347044 225684 347096 225690
rect 347044 225626 347096 225632
rect 346860 178560 346912 178566
rect 346860 178502 346912 178508
rect 346768 113280 346820 113286
rect 346768 113222 346820 113228
rect 348436 89690 348464 322662
rect 349068 254176 349120 254182
rect 349068 254118 349120 254124
rect 348424 89684 348476 89690
rect 348424 89626 348476 89632
rect 346492 36372 346544 36378
rect 346492 36314 346544 36320
rect 346308 36100 346360 36106
rect 346308 36042 346360 36048
rect 344652 12436 344704 12442
rect 344652 12378 344704 12384
rect 343916 8560 343968 8566
rect 343916 8502 343968 8508
rect 342444 5296 342496 5302
rect 342444 5238 342496 5244
rect 339960 5024 340012 5030
rect 339960 4966 340012 4972
rect 349080 3670 349108 254118
rect 349816 195430 349844 505106
rect 351472 496262 351500 525166
rect 351748 524754 351776 525166
rect 351736 524748 351788 524754
rect 351736 524690 351788 524696
rect 351460 496256 351512 496262
rect 351460 496198 351512 496204
rect 351184 306400 351236 306406
rect 351184 306342 351236 306348
rect 349804 195424 349856 195430
rect 349804 195366 349856 195372
rect 349804 187740 349856 187746
rect 349804 187682 349856 187688
rect 349816 4486 349844 187682
rect 351196 13802 351224 306342
rect 351932 119338 351960 619534
rect 352760 619426 352788 619534
rect 352902 619520 353014 620960
rect 356030 619520 356142 620960
rect 358974 619520 359086 620960
rect 362102 619520 362214 620960
rect 365046 619520 365158 620960
rect 367112 619534 367876 619562
rect 352944 619426 352972 619520
rect 352760 619398 352972 619426
rect 356072 616622 356100 619520
rect 356060 616616 356112 616622
rect 356060 616558 356112 616564
rect 363604 616548 363656 616554
rect 363604 616490 363656 616496
rect 359464 616140 359516 616146
rect 359464 616082 359516 616088
rect 355600 529032 355652 529038
rect 355600 528974 355652 528980
rect 355508 528896 355560 528902
rect 355508 528838 355560 528844
rect 353944 527944 353996 527950
rect 353944 527886 353996 527892
rect 353956 385014 353984 527886
rect 353944 385008 353996 385014
rect 353944 384950 353996 384956
rect 355520 119406 355548 528838
rect 355612 365158 355640 528974
rect 358084 460964 358136 460970
rect 358084 460906 358136 460912
rect 356704 457632 356756 457638
rect 356704 457574 356756 457580
rect 355600 365152 355652 365158
rect 355600 365094 355652 365100
rect 355508 119400 355560 119406
rect 355508 119342 355560 119348
rect 351920 119332 351972 119338
rect 351920 119274 351972 119280
rect 356716 23458 356744 457574
rect 357348 148232 357400 148238
rect 357348 148174 357400 148180
rect 356796 128648 356848 128654
rect 356796 128590 356848 128596
rect 356704 23452 356756 23458
rect 356704 23394 356756 23400
rect 351184 13796 351236 13802
rect 351184 13738 351236 13744
rect 349804 4480 349856 4486
rect 349804 4422 349856 4428
rect 338028 3664 338080 3670
rect 338028 3606 338080 3612
rect 348332 3664 348384 3670
rect 348332 3606 348384 3612
rect 349068 3664 349120 3670
rect 349068 3606 349120 3612
rect 342260 3256 342312 3262
rect 342260 3198 342312 3204
rect 333520 3052 333572 3058
rect 333520 2994 333572 3000
rect 342272 480 342300 3198
rect 348344 480 348372 3606
rect 356808 3058 356836 128590
rect 356796 3052 356848 3058
rect 356796 2994 356848 3000
rect 354220 2916 354272 2922
rect 354220 2858 354272 2864
rect 354232 480 354260 2858
rect 357360 2854 357388 148174
rect 358096 106350 358124 460906
rect 358084 106344 358136 106350
rect 358084 106286 358136 106292
rect 359476 70446 359504 616082
rect 363512 545148 363564 545154
rect 363512 545090 363564 545096
rect 361488 533996 361540 534002
rect 361488 533938 361540 533944
rect 360568 475788 360620 475794
rect 360568 475730 360620 475736
rect 360384 394732 360436 394738
rect 360384 394674 360436 394680
rect 360396 366450 360424 394674
rect 360580 366586 360608 475730
rect 360568 366580 360620 366586
rect 360568 366522 360620 366528
rect 360384 366444 360436 366450
rect 360384 366386 360436 366392
rect 360200 366376 360252 366382
rect 360200 366318 360252 366324
rect 359464 70440 359516 70446
rect 359464 70382 359516 70388
rect 360108 66496 360160 66502
rect 360108 66438 360160 66444
rect 360120 9246 360148 66438
rect 360212 25158 360240 366318
rect 360396 339250 360424 366386
rect 361500 359922 361528 533938
rect 361488 359916 361540 359922
rect 361488 359858 361540 359864
rect 361672 359712 361724 359718
rect 361672 359654 361724 359660
rect 361580 356040 361632 356046
rect 361580 355982 361632 355988
rect 360384 339244 360436 339250
rect 360384 339186 360436 339192
rect 360844 325780 360896 325786
rect 360844 325722 360896 325728
rect 360856 124710 360884 325722
rect 361592 250034 361620 355982
rect 361580 250028 361632 250034
rect 361580 249970 361632 249976
rect 361684 220182 361712 359654
rect 363524 331226 363552 545090
rect 363512 331220 363564 331226
rect 363512 331162 363564 331168
rect 362224 222216 362276 222222
rect 362224 222158 362276 222164
rect 361672 220176 361724 220182
rect 361672 220118 361724 220124
rect 361488 142792 361540 142798
rect 361488 142734 361540 142740
rect 360844 124704 360896 124710
rect 360844 124646 360896 124652
rect 360200 25152 360252 25158
rect 360200 25094 360252 25100
rect 360108 9240 360160 9246
rect 360108 9182 360160 9188
rect 361500 3670 361528 142734
rect 362236 72690 362264 222158
rect 363616 126478 363644 616490
rect 364248 614984 364300 614990
rect 364248 614926 364300 614932
rect 363604 126472 363656 126478
rect 363604 126414 363656 126420
rect 362224 72684 362276 72690
rect 362224 72626 362276 72632
rect 360292 3664 360344 3670
rect 360292 3606 360344 3612
rect 361488 3664 361540 3670
rect 361488 3606 361540 3612
rect 363420 3664 363472 3670
rect 363420 3606 363472 3612
rect 357348 2848 357400 2854
rect 357348 2790 357400 2796
rect 360304 480 360332 3606
rect 363432 480 363460 3606
rect 364260 2922 364288 614926
rect 367008 491632 367060 491638
rect 367008 491574 367060 491580
rect 366732 375488 366784 375494
rect 366732 375430 366784 375436
rect 366364 351688 366416 351694
rect 366364 351630 366416 351636
rect 365812 334688 365864 334694
rect 365812 334630 365864 334636
rect 365824 3670 365852 334630
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 366376 3262 366404 351630
rect 366744 123282 366772 375430
rect 366824 371680 366876 371686
rect 366824 371622 366876 371628
rect 366836 123418 366864 371622
rect 366824 123412 366876 123418
rect 366824 123354 366876 123360
rect 366732 123276 366784 123282
rect 366732 123218 366784 123224
rect 366744 108526 366772 123218
rect 367020 123214 367048 491574
rect 367112 292942 367140 619534
rect 367848 619426 367876 619534
rect 367990 619520 368102 620960
rect 371118 619520 371230 620960
rect 374062 619520 374174 620960
rect 377190 619520 377302 620960
rect 379532 619534 380020 619562
rect 368032 619426 368060 619520
rect 367848 619398 368060 619426
rect 371160 617574 371188 619520
rect 369860 617568 369912 617574
rect 369860 617510 369912 617516
rect 371148 617568 371200 617574
rect 371148 617510 371200 617516
rect 367744 541544 367796 541550
rect 367744 541486 367796 541492
rect 367756 387122 367784 541486
rect 369124 500608 369176 500614
rect 369124 500550 369176 500556
rect 367744 387116 367796 387122
rect 367744 387058 367796 387064
rect 368388 387048 368440 387054
rect 368388 386990 368440 386996
rect 367560 386980 367612 386986
rect 367560 386922 367612 386928
rect 367100 292936 367152 292942
rect 367100 292878 367152 292884
rect 367572 282198 367600 386922
rect 368020 386912 368072 386918
rect 368020 386854 368072 386860
rect 367560 282192 367612 282198
rect 367560 282134 367612 282140
rect 367284 266824 367336 266830
rect 367284 266766 367336 266772
rect 367468 266824 367520 266830
rect 367468 266766 367520 266772
rect 367296 223378 367324 266766
rect 367284 223372 367336 223378
rect 367284 223314 367336 223320
rect 367008 123208 367060 123214
rect 367008 123150 367060 123156
rect 367100 123208 367152 123214
rect 367100 123150 367152 123156
rect 366732 108520 366784 108526
rect 366732 108462 366784 108468
rect 367020 50318 367048 123150
rect 367112 111314 367140 123150
rect 367100 111308 367152 111314
rect 367100 111250 367152 111256
rect 367480 72486 367508 266766
rect 368032 108458 368060 386854
rect 368020 108452 368072 108458
rect 368020 108394 368072 108400
rect 368400 105466 368428 386990
rect 368388 105460 368440 105466
rect 368388 105402 368440 105408
rect 368400 105126 368428 105402
rect 368388 105120 368440 105126
rect 368388 105062 368440 105068
rect 369136 84658 369164 500550
rect 369216 282056 369268 282062
rect 369216 281998 369268 282004
rect 369124 84652 369176 84658
rect 369124 84594 369176 84600
rect 367468 72480 367520 72486
rect 367468 72422 367520 72428
rect 367008 50312 367060 50318
rect 367008 50254 367060 50260
rect 369228 45558 369256 281998
rect 369308 133000 369360 133006
rect 369308 132942 369360 132948
rect 369216 45552 369268 45558
rect 369216 45494 369268 45500
rect 368480 36712 368532 36718
rect 368480 36654 368532 36660
rect 368492 16574 368520 36654
rect 368492 16546 369072 16574
rect 366364 3256 366416 3262
rect 366364 3198 366416 3204
rect 364248 2916 364300 2922
rect 364248 2858 364300 2864
rect 369044 490 369072 16546
rect 369320 3670 369348 132942
rect 369872 117774 369900 617510
rect 371792 616412 371844 616418
rect 371792 616354 371844 616360
rect 371240 387116 371292 387122
rect 371240 387058 371292 387064
rect 371148 256080 371200 256086
rect 371148 256022 371200 256028
rect 371160 216986 371188 256022
rect 371148 216980 371200 216986
rect 371148 216922 371200 216928
rect 371160 216782 371188 216922
rect 371148 216776 371200 216782
rect 371148 216718 371200 216724
rect 369860 117768 369912 117774
rect 369860 117710 369912 117716
rect 370504 112396 370556 112402
rect 370504 112338 370556 112344
rect 370516 72622 370544 112338
rect 370504 72616 370556 72622
rect 370504 72558 370556 72564
rect 371252 4146 371280 387058
rect 371424 256012 371476 256018
rect 371424 255954 371476 255960
rect 371436 216782 371464 255954
rect 371424 216776 371476 216782
rect 371424 216718 371476 216724
rect 371804 34746 371832 616354
rect 374104 605834 374132 619520
rect 374012 605806 374132 605834
rect 372712 580576 372764 580582
rect 372712 580518 372764 580524
rect 372620 238536 372672 238542
rect 372620 238478 372672 238484
rect 372632 237454 372660 238478
rect 372620 237448 372672 237454
rect 372620 237390 372672 237396
rect 372632 105330 372660 237390
rect 372620 105324 372672 105330
rect 372620 105266 372672 105272
rect 372724 59634 372752 580518
rect 373816 507204 373868 507210
rect 373816 507146 373868 507152
rect 373080 271380 373132 271386
rect 373080 271322 373132 271328
rect 373092 271182 373120 271322
rect 373080 271176 373132 271182
rect 373080 271118 373132 271124
rect 373092 238542 373120 271118
rect 373828 270842 373856 507146
rect 373816 270836 373868 270842
rect 373816 270778 373868 270784
rect 373080 238536 373132 238542
rect 373080 238478 373132 238484
rect 374012 220561 374040 605806
rect 376484 569288 376536 569294
rect 376484 569230 376536 569236
rect 376208 553444 376260 553450
rect 376208 553386 376260 553392
rect 375656 527264 375708 527270
rect 375656 527206 375708 527212
rect 375668 410446 375696 527206
rect 376220 441998 376248 553386
rect 376208 441992 376260 441998
rect 376208 441934 376260 441940
rect 376116 441856 376168 441862
rect 376116 441798 376168 441804
rect 375380 410440 375432 410446
rect 375380 410382 375432 410388
rect 375656 410440 375708 410446
rect 375656 410382 375708 410388
rect 373998 220552 374054 220561
rect 373998 220487 374054 220496
rect 372712 59628 372764 59634
rect 372712 59570 372764 59576
rect 373172 36168 373224 36174
rect 373172 36110 373224 36116
rect 371792 34740 371844 34746
rect 371792 34682 371844 34688
rect 371804 10470 371832 34682
rect 373184 34610 373212 36110
rect 372896 34604 372948 34610
rect 372896 34546 372948 34552
rect 373172 34604 373224 34610
rect 373172 34546 373224 34552
rect 372908 26234 372936 34546
rect 372908 26206 373028 26234
rect 371792 10464 371844 10470
rect 371792 10406 371844 10412
rect 373000 9042 373028 26206
rect 372988 9036 373040 9042
rect 372988 8978 373040 8984
rect 371240 4140 371292 4146
rect 371240 4082 371292 4088
rect 372436 4140 372488 4146
rect 372436 4082 372488 4088
rect 369308 3664 369360 3670
rect 369308 3606 369360 3612
rect 369320 598 369532 626
rect 369320 490 369348 598
rect 320886 -960 320998 480
rect 324014 -960 324126 480
rect 326958 -960 327070 480
rect 330086 -960 330198 480
rect 333030 -960 333142 480
rect 336158 -960 336270 480
rect 339102 -960 339214 480
rect 342230 -960 342342 480
rect 345174 -960 345286 480
rect 348302 -960 348414 480
rect 351246 -960 351358 480
rect 354190 -960 354302 480
rect 357318 -960 357430 480
rect 360262 -960 360374 480
rect 363390 -960 363502 480
rect 366334 -960 366446 480
rect 369044 462 369348 490
rect 369504 480 369532 598
rect 372448 480 372476 4082
rect 375392 3641 375420 410382
rect 376128 399566 376156 441798
rect 375472 399560 375524 399566
rect 375472 399502 375524 399508
rect 376116 399560 376168 399566
rect 376116 399502 376168 399508
rect 375484 271386 375512 399502
rect 375472 271380 375524 271386
rect 375472 271322 375524 271328
rect 376220 67590 376248 441934
rect 376208 67584 376260 67590
rect 376208 67526 376260 67532
rect 376024 27464 376076 27470
rect 376024 27406 376076 27412
rect 375378 3632 375434 3641
rect 376036 3602 376064 27406
rect 376496 5098 376524 569230
rect 379244 547392 379296 547398
rect 379244 547334 379296 547340
rect 379256 541618 379284 547334
rect 379244 541612 379296 541618
rect 379244 541554 379296 541560
rect 378784 491700 378836 491706
rect 378784 491642 378836 491648
rect 378796 161974 378824 491642
rect 379532 223446 379560 619534
rect 379992 619426 380020 619534
rect 380134 619520 380246 620960
rect 382292 619534 383148 619562
rect 380176 619426 380204 619520
rect 379992 619398 380204 619426
rect 380624 547528 380676 547534
rect 380624 547470 380676 547476
rect 380636 527474 380664 547470
rect 380624 527468 380676 527474
rect 380624 527410 380676 527416
rect 380636 527202 380664 527410
rect 380624 527196 380676 527202
rect 380624 527138 380676 527144
rect 380716 495916 380768 495922
rect 380716 495858 380768 495864
rect 380624 395276 380676 395282
rect 380624 395218 380676 395224
rect 379520 223440 379572 223446
rect 379520 223382 379572 223388
rect 380636 162042 380664 395218
rect 380728 395214 380756 495858
rect 380716 395208 380768 395214
rect 380716 395150 380768 395156
rect 380900 395072 380952 395078
rect 380900 395014 380952 395020
rect 380912 308650 380940 395014
rect 381452 329452 381504 329458
rect 381452 329394 381504 329400
rect 381464 329050 381492 329394
rect 381452 329044 381504 329050
rect 381452 328986 381504 328992
rect 380900 308644 380952 308650
rect 380900 308586 380952 308592
rect 381464 255270 381492 328986
rect 381452 255264 381504 255270
rect 381452 255206 381504 255212
rect 382292 223174 382320 619534
rect 383120 619426 383148 619534
rect 383262 619520 383374 620960
rect 386206 619520 386318 620960
rect 389334 619520 389446 620960
rect 392278 619520 392390 620960
rect 395406 619520 395518 620960
rect 398350 619520 398462 620960
rect 401478 619520 401590 620960
rect 404422 619520 404534 620960
rect 407366 619520 407478 620960
rect 410494 619520 410606 620960
rect 412652 619534 413324 619562
rect 383304 619426 383332 619520
rect 383120 619398 383332 619426
rect 382556 616616 382608 616622
rect 382556 616558 382608 616564
rect 382568 482458 382596 616558
rect 386420 609544 386472 609550
rect 386420 609486 386472 609492
rect 383660 527196 383712 527202
rect 383660 527138 383712 527144
rect 383672 518894 383700 527138
rect 383672 518866 383976 518894
rect 383948 507686 383976 518866
rect 383936 507680 383988 507686
rect 383936 507622 383988 507628
rect 383844 504416 383896 504422
rect 383844 504358 383896 504364
rect 382556 482452 382608 482458
rect 382556 482394 382608 482400
rect 382280 223168 382332 223174
rect 382280 223110 382332 223116
rect 381084 222284 381136 222290
rect 381084 222226 381136 222232
rect 381096 162042 381124 222226
rect 380624 162036 380676 162042
rect 380624 161978 380676 161984
rect 381084 162036 381136 162042
rect 381084 161978 381136 161984
rect 378784 161968 378836 161974
rect 378784 161910 378836 161916
rect 380164 161832 380216 161838
rect 380164 161774 380216 161780
rect 382188 161832 382240 161838
rect 382188 161774 382240 161780
rect 380176 112470 380204 161774
rect 380164 112464 380216 112470
rect 380164 112406 380216 112412
rect 382200 85814 382228 161774
rect 382188 85808 382240 85814
rect 382188 85750 382240 85756
rect 378968 72616 379020 72622
rect 378968 72558 379020 72564
rect 378980 72486 379008 72558
rect 382200 72486 382228 85750
rect 378968 72480 379020 72486
rect 378968 72422 379020 72428
rect 382188 72480 382240 72486
rect 382188 72422 382240 72428
rect 376668 67584 376720 67590
rect 376668 67526 376720 67532
rect 376680 66638 376708 67526
rect 376668 66632 376720 66638
rect 376668 66574 376720 66580
rect 378980 44946 379008 72422
rect 378968 44940 379020 44946
rect 378968 44882 379020 44888
rect 382568 9314 382596 482394
rect 383752 482112 383804 482118
rect 383752 482054 383804 482060
rect 383764 10334 383792 482054
rect 383856 448390 383884 504358
rect 383948 482322 383976 507622
rect 384028 504620 384080 504626
rect 384028 504562 384080 504568
rect 383936 482316 383988 482322
rect 383936 482258 383988 482264
rect 383844 448384 383896 448390
rect 383844 448326 383896 448332
rect 383948 446894 383976 482258
rect 384040 470694 384068 504562
rect 384304 491972 384356 491978
rect 384304 491914 384356 491920
rect 384028 470688 384080 470694
rect 384028 470630 384080 470636
rect 383936 446888 383988 446894
rect 383936 446830 383988 446836
rect 384316 124778 384344 491914
rect 385132 423428 385184 423434
rect 385132 423370 385184 423376
rect 385144 338162 385172 423370
rect 385132 338156 385184 338162
rect 385132 338098 385184 338104
rect 385224 338156 385276 338162
rect 385224 338098 385276 338104
rect 385236 334354 385264 338098
rect 385224 334348 385276 334354
rect 385224 334290 385276 334296
rect 385224 325100 385276 325106
rect 385224 325042 385276 325048
rect 385040 325032 385092 325038
rect 385040 324974 385092 324980
rect 385052 161906 385080 324974
rect 385236 161906 385264 325042
rect 385040 161900 385092 161906
rect 385040 161842 385092 161848
rect 385224 161900 385276 161906
rect 385224 161842 385276 161848
rect 385592 161900 385644 161906
rect 385592 161842 385644 161848
rect 385776 161900 385828 161906
rect 385776 161842 385828 161848
rect 384304 124772 384356 124778
rect 384304 124714 384356 124720
rect 384304 117972 384356 117978
rect 384304 117914 384356 117920
rect 384316 37874 384344 117914
rect 385236 50182 385264 161842
rect 385604 121922 385632 161842
rect 385592 121916 385644 121922
rect 385592 121858 385644 121864
rect 385788 119474 385816 161842
rect 385776 119468 385828 119474
rect 385776 119410 385828 119416
rect 385224 50176 385276 50182
rect 385224 50118 385276 50124
rect 384304 37868 384356 37874
rect 384304 37810 384356 37816
rect 386432 16574 386460 609486
rect 389376 605834 389404 619520
rect 392320 616690 392348 619520
rect 392308 616684 392360 616690
rect 392308 616626 392360 616632
rect 393228 616684 393280 616690
rect 393228 616626 393280 616632
rect 389824 616412 389876 616418
rect 389824 616354 389876 616360
rect 389192 605806 389404 605834
rect 388444 541000 388496 541006
rect 388444 540942 388496 540948
rect 388456 100774 388484 540942
rect 389192 411942 389220 605806
rect 389180 411936 389232 411942
rect 389180 411878 389232 411884
rect 389364 143200 389416 143206
rect 389364 143142 389416 143148
rect 388444 100768 388496 100774
rect 388444 100710 388496 100716
rect 386432 16546 387288 16574
rect 383752 10328 383804 10334
rect 383752 10270 383804 10276
rect 382556 9308 382608 9314
rect 382556 9250 382608 9256
rect 384580 7608 384632 7614
rect 384580 7550 384632 7556
rect 376484 5092 376536 5098
rect 376484 5034 376536 5040
rect 375378 3567 375434 3576
rect 376024 3596 376076 3602
rect 376024 3538 376076 3544
rect 375564 2984 375616 2990
rect 375564 2926 375616 2932
rect 375576 480 375604 2926
rect 384592 480 384620 7550
rect 387260 490 387288 16546
rect 389376 3738 389404 143142
rect 389836 7886 389864 616354
rect 393240 339726 393268 616626
rect 395344 616140 395396 616146
rect 395344 616082 395396 616088
rect 393228 339720 393280 339726
rect 393228 339662 393280 339668
rect 390928 334280 390980 334286
rect 390928 334222 390980 334228
rect 390940 35290 390968 334222
rect 392124 295520 392176 295526
rect 392124 295462 392176 295468
rect 392136 35894 392164 295462
rect 393320 291372 393372 291378
rect 393320 291314 393372 291320
rect 393332 111926 393360 291314
rect 393320 111920 393372 111926
rect 393320 111862 393372 111868
rect 392044 35866 392164 35894
rect 390928 35284 390980 35290
rect 390928 35226 390980 35232
rect 392044 35086 392072 35866
rect 392032 35080 392084 35086
rect 392032 35022 392084 35028
rect 393332 16574 393360 111862
rect 395356 37670 395384 616082
rect 396724 578944 396776 578950
rect 396724 578886 396776 578892
rect 396632 254856 396684 254862
rect 396632 254798 396684 254804
rect 396644 99278 396672 254798
rect 396736 112810 396764 578886
rect 400036 398472 400088 398478
rect 400036 398414 400088 398420
rect 398104 396296 398156 396302
rect 398104 396238 398156 396244
rect 396724 112804 396776 112810
rect 396724 112746 396776 112752
rect 396632 99272 396684 99278
rect 396632 99214 396684 99220
rect 398116 59226 398144 396238
rect 400048 322930 400076 398414
rect 401140 333056 401192 333062
rect 401140 332998 401192 333004
rect 400036 322924 400088 322930
rect 400036 322866 400088 322872
rect 399484 218068 399536 218074
rect 399484 218010 399536 218016
rect 398104 59220 398156 59226
rect 398104 59162 398156 59168
rect 395344 37664 395396 37670
rect 395344 37606 395396 37612
rect 399496 32026 399524 218010
rect 401152 54534 401180 332998
rect 401520 320210 401548 619520
rect 404464 616078 404492 619520
rect 404452 616072 404504 616078
rect 404452 616014 404504 616020
rect 402428 611720 402480 611726
rect 402428 611662 402480 611668
rect 402440 414254 402468 611662
rect 405924 583432 405976 583438
rect 405924 583374 405976 583380
rect 403440 578944 403492 578950
rect 403440 578886 403492 578892
rect 403452 557394 403480 578886
rect 403440 557388 403492 557394
rect 403440 557330 403492 557336
rect 403348 557184 403400 557190
rect 403348 557126 403400 557132
rect 402980 534336 403032 534342
rect 402980 534278 403032 534284
rect 402428 414248 402480 414254
rect 402428 414190 402480 414196
rect 402440 356046 402468 414190
rect 402992 360398 403020 534278
rect 402796 360392 402848 360398
rect 402796 360334 402848 360340
rect 402980 360392 403032 360398
rect 402980 360334 403032 360340
rect 402428 356040 402480 356046
rect 402428 355982 402480 355988
rect 401508 320204 401560 320210
rect 401508 320146 401560 320152
rect 402808 273970 402836 360334
rect 402796 273964 402848 273970
rect 402796 273906 402848 273912
rect 402992 262478 403020 360334
rect 402980 262472 403032 262478
rect 402980 262414 403032 262420
rect 403360 112538 403388 557126
rect 403452 556238 403480 557330
rect 403440 556232 403492 556238
rect 403440 556174 403492 556180
rect 404268 534744 404320 534750
rect 404268 534686 404320 534692
rect 404280 534342 404308 534686
rect 404268 534336 404320 534342
rect 404268 534278 404320 534284
rect 405832 514344 405884 514350
rect 405832 514286 405884 514292
rect 405372 514208 405424 514214
rect 405372 514150 405424 514156
rect 403808 414112 403860 414118
rect 403808 414054 403860 414060
rect 403820 384334 403848 414054
rect 403808 384328 403860 384334
rect 403808 384270 403860 384276
rect 405004 375080 405056 375086
rect 405004 375022 405056 375028
rect 403348 112532 403400 112538
rect 403348 112474 403400 112480
rect 401232 59560 401284 59566
rect 401232 59502 401284 59508
rect 401244 54670 401272 59502
rect 401232 54664 401284 54670
rect 401232 54606 401284 54612
rect 401140 54528 401192 54534
rect 401140 54470 401192 54476
rect 399484 32020 399536 32026
rect 399484 31962 399536 31968
rect 393332 16546 393636 16574
rect 389824 7880 389876 7886
rect 389824 7822 389876 7828
rect 389364 3732 389416 3738
rect 389364 3674 389416 3680
rect 390652 2848 390704 2854
rect 390652 2790 390704 2796
rect 387536 598 387748 626
rect 387536 490 387564 598
rect 369462 -960 369574 480
rect 372406 -960 372518 480
rect 375534 -960 375646 480
rect 378478 -960 378590 480
rect 381606 -960 381718 480
rect 384550 -960 384662 480
rect 387260 462 387564 490
rect 387720 480 387748 598
rect 390664 480 390692 2790
rect 393608 480 393636 16546
rect 401244 9110 401272 54606
rect 401232 9104 401284 9110
rect 401232 9046 401284 9052
rect 405016 8226 405044 375022
rect 405384 8634 405412 514150
rect 405740 113008 405792 113014
rect 405740 112950 405792 112956
rect 405372 8628 405424 8634
rect 405372 8570 405424 8576
rect 405004 8220 405056 8226
rect 405004 8162 405056 8168
rect 405752 480 405780 112950
rect 405844 112878 405872 514286
rect 405936 197334 405964 583374
rect 406016 556232 406068 556238
rect 406016 556174 406068 556180
rect 406028 514350 406056 556174
rect 406016 514344 406068 514350
rect 406016 514286 406068 514292
rect 409604 514344 409656 514350
rect 409604 514286 409656 514292
rect 406568 504620 406620 504626
rect 406568 504562 406620 504568
rect 406580 503742 406608 504562
rect 406568 503736 406620 503742
rect 406568 503678 406620 503684
rect 406292 280492 406344 280498
rect 406292 280434 406344 280440
rect 405924 197328 405976 197334
rect 405924 197270 405976 197276
rect 405832 112872 405884 112878
rect 405832 112814 405884 112820
rect 406304 59770 406332 280434
rect 406384 271108 406436 271114
rect 406384 271050 406436 271056
rect 406396 179790 406424 271050
rect 406384 179784 406436 179790
rect 406384 179726 406436 179732
rect 406396 78538 406424 179726
rect 406384 78532 406436 78538
rect 406384 78474 406436 78480
rect 406580 64874 406608 503678
rect 407396 387524 407448 387530
rect 407396 387466 407448 387472
rect 407408 179654 407436 387466
rect 409420 375148 409472 375154
rect 409420 375090 409472 375096
rect 409052 374944 409104 374950
rect 409052 374886 409104 374892
rect 407396 179648 407448 179654
rect 407396 179590 407448 179596
rect 407408 178226 407436 179590
rect 407396 178220 407448 178226
rect 407396 178162 407448 178168
rect 409064 110702 409092 374886
rect 409432 118046 409460 375090
rect 409616 375086 409644 514286
rect 410524 513800 410576 513806
rect 410524 513742 410576 513748
rect 409604 375080 409656 375086
rect 409604 375022 409656 375028
rect 409420 118040 409472 118046
rect 409420 117982 409472 117988
rect 409052 110696 409104 110702
rect 409052 110638 409104 110644
rect 406488 64846 406608 64874
rect 406292 59764 406344 59770
rect 406292 59706 406344 59712
rect 406304 59634 406332 59706
rect 406488 59634 406516 64846
rect 406292 59628 406344 59634
rect 406292 59570 406344 59576
rect 406476 59628 406528 59634
rect 406476 59570 406528 59576
rect 410536 35902 410564 513742
rect 412088 439884 412140 439890
rect 412088 439826 412140 439832
rect 412100 428262 412128 439826
rect 412272 439748 412324 439754
rect 412272 439690 412324 439696
rect 412284 428466 412312 439690
rect 412272 428460 412324 428466
rect 412272 428402 412324 428408
rect 412364 428460 412416 428466
rect 412364 428402 412416 428408
rect 412088 428256 412140 428262
rect 412088 428198 412140 428204
rect 412100 120086 412128 428198
rect 412284 387190 412312 428402
rect 412272 387184 412324 387190
rect 412272 387126 412324 387132
rect 412376 312118 412404 428402
rect 412364 312112 412416 312118
rect 412364 312054 412416 312060
rect 412088 120080 412140 120086
rect 412088 120022 412140 120028
rect 412652 118182 412680 619534
rect 413296 619426 413324 619534
rect 413438 619520 413550 620960
rect 416566 619520 416678 620960
rect 419510 619520 419622 620960
rect 422638 619520 422750 620960
rect 425582 619520 425694 620960
rect 428710 619520 428822 620960
rect 430592 619534 431540 619562
rect 413480 619426 413508 619520
rect 413296 619398 413508 619426
rect 416608 616486 416636 619520
rect 428752 616826 428780 619520
rect 428740 616820 428792 616826
rect 428740 616762 428792 616768
rect 416596 616480 416648 616486
rect 416596 616422 416648 616428
rect 425704 616344 425756 616350
rect 425704 616286 425756 616292
rect 419540 610224 419592 610230
rect 419540 610166 419592 610172
rect 419552 590646 419580 610166
rect 419540 590640 419592 590646
rect 419540 590582 419592 590588
rect 419356 590572 419408 590578
rect 419356 590514 419408 590520
rect 416688 586900 416740 586906
rect 416688 586842 416740 586848
rect 416596 544264 416648 544270
rect 416596 544206 416648 544212
rect 412916 489864 412968 489870
rect 412916 489806 412968 489812
rect 412928 482254 412956 489806
rect 414296 489728 414348 489734
rect 414296 489670 414348 489676
rect 412916 482248 412968 482254
rect 412916 482190 412968 482196
rect 414308 400722 414336 489670
rect 414296 400716 414348 400722
rect 414296 400658 414348 400664
rect 414388 384464 414440 384470
rect 414388 384406 414440 384412
rect 414400 296206 414428 384406
rect 414388 296200 414440 296206
rect 414388 296142 414440 296148
rect 414664 252680 414716 252686
rect 414664 252622 414716 252628
rect 412640 118176 412692 118182
rect 412640 118118 412692 118124
rect 410524 35896 410576 35902
rect 410524 35838 410576 35844
rect 414676 13870 414704 252622
rect 416136 236360 416188 236366
rect 416136 236302 416188 236308
rect 414848 161696 414900 161702
rect 414848 161638 414900 161644
rect 414664 13864 414716 13870
rect 414664 13806 414716 13812
rect 414860 4010 414888 161638
rect 416148 140622 416176 236302
rect 416136 140616 416188 140622
rect 416136 140558 416188 140564
rect 416412 140548 416464 140554
rect 416412 140490 416464 140496
rect 416424 111450 416452 140490
rect 416412 111444 416464 111450
rect 416412 111386 416464 111392
rect 416608 108322 416636 544206
rect 416596 108316 416648 108322
rect 416596 108258 416648 108264
rect 416700 31482 416728 586842
rect 417884 570784 417936 570790
rect 417884 570726 417936 570732
rect 417792 527808 417844 527814
rect 417792 527750 417844 527756
rect 417804 487286 417832 527750
rect 417896 487286 417924 570726
rect 417976 529032 418028 529038
rect 417976 528974 418028 528980
rect 417792 487280 417844 487286
rect 417792 487222 417844 487228
rect 417884 487280 417936 487286
rect 417884 487222 417936 487228
rect 417804 329798 417832 487222
rect 417516 329792 417568 329798
rect 417516 329734 417568 329740
rect 417792 329792 417844 329798
rect 417792 329734 417844 329740
rect 417528 329322 417556 329734
rect 417896 329594 417924 487222
rect 417988 487218 418016 528974
rect 417976 487212 418028 487218
rect 417976 487154 418028 487160
rect 419368 448526 419396 590514
rect 419632 590368 419684 590374
rect 419632 590310 419684 590316
rect 419356 448520 419408 448526
rect 419356 448462 419408 448468
rect 418804 439816 418856 439822
rect 418804 439758 418856 439764
rect 417884 329588 417936 329594
rect 417884 329530 417936 329536
rect 417516 329316 417568 329322
rect 417516 329258 417568 329264
rect 418712 230784 418764 230790
rect 418712 230726 418764 230732
rect 417516 152040 417568 152046
rect 417516 151982 417568 151988
rect 417424 140480 417476 140486
rect 417424 140422 417476 140428
rect 417436 111382 417464 140422
rect 417424 111376 417476 111382
rect 417424 111318 417476 111324
rect 416872 35080 416924 35086
rect 416872 35022 416924 35028
rect 416688 31476 416740 31482
rect 416688 31418 416740 31424
rect 416884 31414 416912 35022
rect 417528 31482 417556 151982
rect 418160 143540 418212 143546
rect 418160 143482 418212 143488
rect 418172 142866 418200 143482
rect 418160 142860 418212 142866
rect 418160 142802 418212 142808
rect 418724 112742 418752 230726
rect 418816 143546 418844 439758
rect 418988 439680 419040 439686
rect 418988 439622 419040 439628
rect 418804 143540 418856 143546
rect 418804 143482 418856 143488
rect 418712 112736 418764 112742
rect 418712 112678 418764 112684
rect 419000 110770 419028 439622
rect 419080 375080 419132 375086
rect 419080 375022 419132 375028
rect 419092 230994 419120 375022
rect 419080 230988 419132 230994
rect 419080 230930 419132 230936
rect 419092 161906 419120 230930
rect 419540 175636 419592 175642
rect 419540 175578 419592 175584
rect 419080 161900 419132 161906
rect 419080 161842 419132 161848
rect 418988 110764 419040 110770
rect 418988 110706 419040 110712
rect 419552 107982 419580 175578
rect 419644 111722 419672 590310
rect 423588 576904 423640 576910
rect 423588 576846 423640 576852
rect 422944 572076 422996 572082
rect 422944 572018 422996 572024
rect 421012 500880 421064 500886
rect 421012 500822 421064 500828
rect 420736 500812 420788 500818
rect 420736 500754 420788 500760
rect 420552 500676 420604 500682
rect 420552 500618 420604 500624
rect 420644 500676 420696 500682
rect 420644 500618 420696 500624
rect 420564 485518 420592 500618
rect 420552 485512 420604 485518
rect 420552 485454 420604 485460
rect 420656 435130 420684 500618
rect 420748 485586 420776 500754
rect 420920 500744 420972 500750
rect 420920 500686 420972 500692
rect 420736 485580 420788 485586
rect 420736 485522 420788 485528
rect 420644 435124 420696 435130
rect 420644 435066 420696 435072
rect 420932 346662 420960 500686
rect 421024 485382 421052 500822
rect 422024 487212 422076 487218
rect 422024 487154 422076 487160
rect 421012 485376 421064 485382
rect 421012 485318 421064 485324
rect 420920 346656 420972 346662
rect 420920 346598 420972 346604
rect 420552 272672 420604 272678
rect 420552 272614 420604 272620
rect 419632 111716 419684 111722
rect 419632 111658 419684 111664
rect 419540 107976 419592 107982
rect 419540 107918 419592 107924
rect 418436 72480 418488 72486
rect 418436 72422 418488 72428
rect 418448 37806 418476 72422
rect 419552 59702 419580 107918
rect 419540 59696 419592 59702
rect 419540 59638 419592 59644
rect 418344 37800 418396 37806
rect 418344 37742 418396 37748
rect 418436 37800 418488 37806
rect 418436 37742 418488 37748
rect 417884 37664 417936 37670
rect 417884 37606 417936 37612
rect 417516 31476 417568 31482
rect 417516 31418 417568 31424
rect 416872 31408 416924 31414
rect 416872 31350 416924 31356
rect 416884 31278 416912 31350
rect 416872 31272 416924 31278
rect 416872 31214 416924 31220
rect 415492 31136 415544 31142
rect 415492 31078 415544 31084
rect 414848 4004 414900 4010
rect 414848 3946 414900 3952
rect 415504 3369 415532 31078
rect 417896 11898 417924 37606
rect 417884 11892 417936 11898
rect 417884 11834 417936 11840
rect 418356 7546 418384 37742
rect 418344 7540 418396 7546
rect 418344 7482 418396 7488
rect 415490 3360 415546 3369
rect 414940 3324 414992 3330
rect 415490 3295 415546 3304
rect 414940 3266 414992 3272
rect 414952 480 414980 3266
rect 420564 3126 420592 272614
rect 422036 57254 422064 487154
rect 422956 61062 422984 572018
rect 423600 496126 423628 576846
rect 423588 496120 423640 496126
rect 423588 496062 423640 496068
rect 423956 489728 424008 489734
rect 423956 489670 424008 489676
rect 423864 443692 423916 443698
rect 423864 443634 423916 443640
rect 423772 400648 423824 400654
rect 423772 400590 423824 400596
rect 423784 327418 423812 400590
rect 423772 327412 423824 327418
rect 423772 327354 423824 327360
rect 423876 324902 423904 443634
rect 423968 327282 423996 489670
rect 424048 443488 424100 443494
rect 424048 443430 424100 443436
rect 423956 327276 424008 327282
rect 423956 327218 424008 327224
rect 423864 324896 423916 324902
rect 423864 324838 423916 324844
rect 424060 162042 424088 443430
rect 424048 162036 424100 162042
rect 424048 161978 424100 161984
rect 425716 152114 425744 616286
rect 426624 507884 426676 507890
rect 426624 507826 426676 507832
rect 426808 507884 426860 507890
rect 426808 507826 426860 507832
rect 425704 152108 425756 152114
rect 425704 152050 425756 152056
rect 426636 126342 426664 507826
rect 426716 399424 426768 399430
rect 426716 399366 426768 399372
rect 426728 308786 426756 399366
rect 426716 308780 426768 308786
rect 426716 308722 426768 308728
rect 426820 222970 426848 507826
rect 426900 507680 426952 507686
rect 426900 507622 426952 507628
rect 426912 337482 426940 507622
rect 429292 491904 429344 491910
rect 429292 491846 429344 491852
rect 426992 361616 427044 361622
rect 426992 361558 427044 361564
rect 426900 337476 426952 337482
rect 426900 337418 426952 337424
rect 427004 308786 427032 361558
rect 426992 308780 427044 308786
rect 426992 308722 427044 308728
rect 427004 296714 427032 308722
rect 426912 296686 427032 296714
rect 426912 279206 426940 296686
rect 426900 279200 426952 279206
rect 426900 279142 426952 279148
rect 426808 222964 426860 222970
rect 426808 222906 426860 222912
rect 428924 216912 428976 216918
rect 428924 216854 428976 216860
rect 426624 126336 426676 126342
rect 426624 126278 426676 126284
rect 428936 124914 428964 216854
rect 429200 152584 429252 152590
rect 429200 152526 429252 152532
rect 429212 124914 429240 152526
rect 429304 124914 429332 491846
rect 430592 223310 430620 619534
rect 431512 619426 431540 619534
rect 431654 619520 431766 620960
rect 434782 619520 434894 620960
rect 437726 619520 437838 620960
rect 440854 619520 440966 620960
rect 443798 619520 443910 620960
rect 446742 619520 446854 620960
rect 449870 619520 449982 620960
rect 452814 619520 452926 620960
rect 455432 619534 455828 619562
rect 431696 619426 431724 619520
rect 431512 619398 431724 619426
rect 443840 616418 443868 619520
rect 443828 616412 443880 616418
rect 443828 616354 443880 616360
rect 438308 616208 438360 616214
rect 438308 616150 438360 616156
rect 435272 610632 435324 610638
rect 435272 610574 435324 610580
rect 434904 610292 434956 610298
rect 434904 610234 434956 610240
rect 434916 551886 434944 610234
rect 435284 551886 435312 610574
rect 435364 590572 435416 590578
rect 435364 590514 435416 590520
rect 435376 551886 435404 590514
rect 434904 551880 434956 551886
rect 434904 551822 434956 551828
rect 435272 551880 435324 551886
rect 435272 551822 435324 551828
rect 435364 551880 435416 551886
rect 435364 551822 435416 551828
rect 434720 551744 434772 551750
rect 434720 551686 434772 551692
rect 430764 533792 430816 533798
rect 430764 533734 430816 533740
rect 430776 237454 430804 533734
rect 432512 489864 432564 489870
rect 432512 489806 432564 489812
rect 432524 469878 432552 489806
rect 432512 469872 432564 469878
rect 432512 469814 432564 469820
rect 433984 395072 434036 395078
rect 433984 395014 434036 395020
rect 432604 344072 432656 344078
rect 432604 344014 432656 344020
rect 430948 237584 431000 237590
rect 430948 237526 431000 237532
rect 430960 237454 430988 237526
rect 430764 237448 430816 237454
rect 430764 237390 430816 237396
rect 430948 237448 431000 237454
rect 430948 237390 431000 237396
rect 430580 223304 430632 223310
rect 430580 223246 430632 223252
rect 430960 220726 430988 237390
rect 430948 220720 431000 220726
rect 430948 220662 431000 220668
rect 430960 219434 430988 220662
rect 430592 219406 430988 219434
rect 428924 124908 428976 124914
rect 428924 124850 428976 124856
rect 429200 124908 429252 124914
rect 429200 124850 429252 124856
rect 429292 124908 429344 124914
rect 429292 124850 429344 124856
rect 429844 78668 429896 78674
rect 429844 78610 429896 78616
rect 429856 75546 429884 78610
rect 429844 75540 429896 75546
rect 429844 75482 429896 75488
rect 429660 75336 429712 75342
rect 429660 75278 429712 75284
rect 429672 67590 429700 75278
rect 429660 67584 429712 67590
rect 429660 67526 429712 67532
rect 422944 61056 422996 61062
rect 422944 60998 422996 61004
rect 422024 57248 422076 57254
rect 422024 57190 422076 57196
rect 430592 46034 430620 219406
rect 432616 93838 432644 344014
rect 432604 93832 432656 93838
rect 432604 93774 432656 93780
rect 433996 90098 434024 395014
rect 434732 119542 434760 551686
rect 434916 359718 434944 551822
rect 434996 551812 435048 551818
rect 434996 551754 435048 551760
rect 435088 551812 435140 551818
rect 435088 551754 435140 551760
rect 434904 359712 434956 359718
rect 434904 359654 434956 359660
rect 434720 119536 434772 119542
rect 434720 119478 434772 119484
rect 433984 90092 434036 90098
rect 433984 90034 434036 90040
rect 430580 46028 430632 46034
rect 430580 45970 430632 45976
rect 435008 3942 435036 551754
rect 435100 514894 435128 551754
rect 435088 514888 435140 514894
rect 435088 514830 435140 514836
rect 435284 237454 435312 551822
rect 436744 434784 436796 434790
rect 436744 434726 436796 434732
rect 435272 237448 435324 237454
rect 435272 237390 435324 237396
rect 436756 90166 436784 434726
rect 438320 329458 438348 616150
rect 440884 610496 440936 610502
rect 440884 610438 440936 610444
rect 438308 329452 438360 329458
rect 438308 329394 438360 329400
rect 438492 329452 438544 329458
rect 438492 329394 438544 329400
rect 438320 118250 438348 329394
rect 438504 222630 438532 329394
rect 439964 329384 440016 329390
rect 439964 329326 440016 329332
rect 438492 222624 438544 222630
rect 438492 222566 438544 222572
rect 438308 118244 438360 118250
rect 438308 118186 438360 118192
rect 436744 90160 436796 90166
rect 436744 90102 436796 90108
rect 439976 89894 440004 329326
rect 440896 99210 440924 610438
rect 445668 571872 445720 571878
rect 445668 571814 445720 571820
rect 443092 504416 443144 504422
rect 443092 504358 443144 504364
rect 442540 421184 442592 421190
rect 442540 421126 442592 421132
rect 441988 372360 442040 372366
rect 441988 372302 442040 372308
rect 442000 332586 442028 372302
rect 441988 332580 442040 332586
rect 441988 332522 442040 332528
rect 440884 99204 440936 99210
rect 440884 99146 440936 99152
rect 439964 89888 440016 89894
rect 439964 89830 440016 89836
rect 442552 78266 442580 421126
rect 443104 79286 443132 504358
rect 443920 469872 443972 469878
rect 443920 469814 443972 469820
rect 443932 421326 443960 469814
rect 443920 421320 443972 421326
rect 443920 421262 443972 421268
rect 444012 252204 444064 252210
rect 444012 252146 444064 252152
rect 444024 118318 444052 252146
rect 444104 252136 444156 252142
rect 444104 252078 444156 252084
rect 444196 252136 444248 252142
rect 444196 252078 444248 252084
rect 444012 118312 444064 118318
rect 444012 118254 444064 118260
rect 443092 79280 443144 79286
rect 443092 79222 443144 79228
rect 442908 79212 442960 79218
rect 442908 79154 442960 79160
rect 442540 78260 442592 78266
rect 442540 78202 442592 78208
rect 442920 54534 442948 79154
rect 443184 79008 443236 79014
rect 443184 78950 443236 78956
rect 443196 59770 443224 78950
rect 443184 59764 443236 59770
rect 443184 59706 443236 59712
rect 442908 54528 442960 54534
rect 442908 54470 442960 54476
rect 444116 8158 444144 252078
rect 444208 230994 444236 252078
rect 444196 230988 444248 230994
rect 444196 230930 444248 230936
rect 445680 61198 445708 571814
rect 447784 553512 447836 553518
rect 447784 553454 447836 553460
rect 445760 308712 445812 308718
rect 445760 308654 445812 308660
rect 445772 308446 445800 308654
rect 445760 308440 445812 308446
rect 445760 308382 445812 308388
rect 445772 66502 445800 308382
rect 445760 66496 445812 66502
rect 445760 66438 445812 66444
rect 445772 64874 445800 66438
rect 445772 64846 446076 64874
rect 446048 61266 446076 64846
rect 446036 61260 446088 61266
rect 446036 61202 446088 61208
rect 445668 61192 445720 61198
rect 445668 61134 445720 61140
rect 445760 61192 445812 61198
rect 445760 61134 445812 61140
rect 445772 9518 445800 61134
rect 447796 15366 447824 553454
rect 449912 424590 449940 619520
rect 452856 616282 452884 619520
rect 452844 616276 452896 616282
rect 452844 616218 452896 616224
rect 451924 566976 451976 566982
rect 451924 566918 451976 566924
rect 449900 424584 449952 424590
rect 449900 424526 449952 424532
rect 451464 423156 451516 423162
rect 451464 423098 451516 423104
rect 450452 387592 450504 387598
rect 450452 387534 450504 387540
rect 450464 374746 450492 387534
rect 450636 386912 450688 386918
rect 450636 386854 450688 386860
rect 450452 374740 450504 374746
rect 450452 374682 450504 374688
rect 450648 374542 450676 386854
rect 450636 374536 450688 374542
rect 450636 374478 450688 374484
rect 451476 349518 451504 423098
rect 451936 394126 451964 566918
rect 452108 525224 452160 525230
rect 452108 525166 452160 525172
rect 452120 394194 452148 525166
rect 452108 394188 452160 394194
rect 452108 394130 452160 394136
rect 451924 394120 451976 394126
rect 451924 394062 451976 394068
rect 451556 393984 451608 393990
rect 451556 393926 451608 393932
rect 451464 349512 451516 349518
rect 451464 349454 451516 349460
rect 451568 119950 451596 393926
rect 453028 183592 453080 183598
rect 453028 183534 453080 183540
rect 451648 140616 451700 140622
rect 451648 140558 451700 140564
rect 451556 119944 451608 119950
rect 451556 119886 451608 119892
rect 451660 117298 451688 140558
rect 451372 117292 451424 117298
rect 451372 117234 451424 117240
rect 451648 117292 451700 117298
rect 451648 117234 451700 117240
rect 450268 117088 450320 117094
rect 450268 117030 450320 117036
rect 447784 15360 447836 15366
rect 447784 15302 447836 15308
rect 450280 10538 450308 117030
rect 451384 113174 451412 117234
rect 451660 116618 451688 117234
rect 451648 116612 451700 116618
rect 451648 116554 451700 116560
rect 451384 113146 451504 113174
rect 450268 10532 450320 10538
rect 450268 10474 450320 10480
rect 445760 9512 445812 9518
rect 445760 9454 445812 9460
rect 451476 8906 451504 113146
rect 453040 109206 453068 183534
rect 453028 109200 453080 109206
rect 453028 109142 453080 109148
rect 453040 15502 453068 109142
rect 453028 15496 453080 15502
rect 453028 15438 453080 15444
rect 455432 9382 455460 619534
rect 455800 619426 455828 619534
rect 455942 619520 456054 620960
rect 458886 619520 458998 620960
rect 462014 619520 462126 620960
rect 464958 619520 465070 620960
rect 468086 619520 468198 620960
rect 471030 619520 471142 620960
rect 474158 619520 474270 620960
rect 477102 619520 477214 620960
rect 480230 619520 480342 620960
rect 483174 619520 483286 620960
rect 486118 619520 486230 620960
rect 489246 619520 489358 620960
rect 491312 619534 492076 619562
rect 455984 619426 456012 619520
rect 455800 619398 456012 619426
rect 462056 616758 462084 619520
rect 465000 617574 465028 619520
rect 463700 617568 463752 617574
rect 463700 617510 463752 617516
rect 464988 617568 465040 617574
rect 464988 617510 465040 617516
rect 462044 616752 462096 616758
rect 462044 616694 462096 616700
rect 456800 610564 456852 610570
rect 456800 610506 456852 610512
rect 456064 111988 456116 111994
rect 456064 111930 456116 111936
rect 456076 16114 456104 111930
rect 456812 99142 456840 610506
rect 463424 587308 463476 587314
rect 463424 587250 463476 587256
rect 463516 587308 463568 587314
rect 463516 587250 463568 587256
rect 463148 587240 463200 587246
rect 463148 587182 463200 587188
rect 463160 539578 463188 587182
rect 462320 539572 462372 539578
rect 462320 539514 462372 539520
rect 463148 539572 463200 539578
rect 463148 539514 463200 539520
rect 462332 539374 462360 539514
rect 463436 539442 463464 587250
rect 463424 539436 463476 539442
rect 463424 539378 463476 539384
rect 462320 539368 462372 539374
rect 462320 539310 462372 539316
rect 462332 308446 462360 539310
rect 462320 308440 462372 308446
rect 462320 308382 462372 308388
rect 458180 116612 458232 116618
rect 458180 116554 458232 116560
rect 458192 99278 458220 116554
rect 460204 112940 460256 112946
rect 460204 112882 460256 112888
rect 458180 99272 458232 99278
rect 458180 99214 458232 99220
rect 456800 99136 456852 99142
rect 456800 99078 456852 99084
rect 458192 31278 458220 99214
rect 458180 31272 458232 31278
rect 458180 31214 458232 31220
rect 456064 16108 456116 16114
rect 456064 16050 456116 16056
rect 460216 14006 460244 112882
rect 463528 31142 463556 587250
rect 463712 332654 463740 617510
rect 468128 616146 468156 619520
rect 471072 616758 471100 619520
rect 471060 616752 471112 616758
rect 471060 616694 471112 616700
rect 471888 616752 471940 616758
rect 471888 616694 471940 616700
rect 468116 616140 468168 616146
rect 468116 616082 468168 616088
rect 469588 543788 469640 543794
rect 469588 543730 469640 543736
rect 464160 503736 464212 503742
rect 464160 503678 464212 503684
rect 464172 484090 464200 503678
rect 464160 484084 464212 484090
rect 464160 484026 464212 484032
rect 464252 484084 464304 484090
rect 464252 484026 464304 484032
rect 463976 483948 464028 483954
rect 463976 483890 464028 483896
rect 463988 469606 464016 483890
rect 463976 469600 464028 469606
rect 463976 469542 464028 469548
rect 463700 332648 463752 332654
rect 463700 332590 463752 332596
rect 464264 59634 464292 484026
rect 464344 483948 464396 483954
rect 464344 483890 464396 483896
rect 464356 381546 464384 483890
rect 464344 381540 464396 381546
rect 464344 381482 464396 381488
rect 468024 359916 468076 359922
rect 468024 359858 468076 359864
rect 468036 240922 468064 359858
rect 468024 240916 468076 240922
rect 468024 240858 468076 240864
rect 467380 240644 467432 240650
rect 467380 240586 467432 240592
rect 467840 240644 467892 240650
rect 467840 240586 467892 240592
rect 467392 202842 467420 240586
rect 467656 240576 467708 240582
rect 467656 240518 467708 240524
rect 467748 240576 467800 240582
rect 467748 240518 467800 240524
rect 467668 223514 467696 240518
rect 467656 223508 467708 223514
rect 467656 223450 467708 223456
rect 467380 202836 467432 202842
rect 467380 202778 467432 202784
rect 464252 59628 464304 59634
rect 464252 59570 464304 59576
rect 463884 48136 463936 48142
rect 463884 48078 463936 48084
rect 463896 36650 463924 48078
rect 463884 36644 463936 36650
rect 463884 36586 463936 36592
rect 466460 36576 466512 36582
rect 466460 36518 466512 36524
rect 463516 31136 463568 31142
rect 463516 31078 463568 31084
rect 460204 14000 460256 14006
rect 460204 13942 460256 13948
rect 455420 9376 455472 9382
rect 455420 9318 455472 9324
rect 451464 8900 451516 8906
rect 451464 8842 451516 8848
rect 444104 8152 444156 8158
rect 444104 8094 444156 8100
rect 463332 4072 463384 4078
rect 463332 4014 463384 4020
rect 434996 3936 435048 3942
rect 434996 3878 435048 3884
rect 460388 3664 460440 3670
rect 460388 3606 460440 3612
rect 439044 3528 439096 3534
rect 439044 3470 439096 3476
rect 436100 3256 436152 3262
rect 436100 3198 436152 3204
rect 420552 3120 420604 3126
rect 420552 3062 420604 3068
rect 417884 3052 417936 3058
rect 417884 2994 417936 3000
rect 417896 480 417924 2994
rect 421012 2916 421064 2922
rect 421012 2858 421064 2864
rect 421024 480 421052 2858
rect 436112 480 436140 3198
rect 439056 480 439084 3470
rect 445116 3392 445168 3398
rect 445116 3334 445168 3340
rect 445128 480 445156 3334
rect 454316 3188 454368 3194
rect 454316 3130 454368 3136
rect 454328 480 454356 3130
rect 460400 480 460428 3606
rect 463344 480 463372 4014
rect 466472 480 466500 36518
rect 467760 8770 467788 240518
rect 467852 118454 467880 240586
rect 467840 118448 467892 118454
rect 467840 118390 467892 118396
rect 467748 8764 467800 8770
rect 467748 8706 467800 8712
rect 468036 8362 468064 240858
rect 469600 78606 469628 543730
rect 470048 489184 470100 489190
rect 470048 489126 470100 489132
rect 469864 183728 469916 183734
rect 469864 183670 469916 183676
rect 469876 78674 469904 183670
rect 469864 78668 469916 78674
rect 469864 78610 469916 78616
rect 469588 78600 469640 78606
rect 469588 78542 469640 78548
rect 469680 78600 469732 78606
rect 469680 78542 469732 78548
rect 469404 78464 469456 78470
rect 469404 78406 469456 78412
rect 469416 9654 469444 78406
rect 469404 9648 469456 9654
rect 469404 9590 469456 9596
rect 469692 9178 469720 78542
rect 469680 9172 469732 9178
rect 469680 9114 469732 9120
rect 468024 8356 468076 8362
rect 468024 8298 468076 8304
rect 470060 4826 470088 489126
rect 470416 421320 470468 421326
rect 470416 421262 470468 421268
rect 470428 364750 470456 421262
rect 470416 364744 470468 364750
rect 470416 364686 470468 364692
rect 470600 348424 470652 348430
rect 470600 348366 470652 348372
rect 470508 257032 470560 257038
rect 470508 256974 470560 256980
rect 470520 161974 470548 256974
rect 470612 256902 470640 348366
rect 470600 256896 470652 256902
rect 470600 256838 470652 256844
rect 470508 161968 470560 161974
rect 470508 161910 470560 161916
rect 470612 109070 470640 256838
rect 470600 109064 470652 109070
rect 470600 109006 470652 109012
rect 471900 107982 471928 616694
rect 480272 608870 480300 619520
rect 480260 608864 480312 608870
rect 480260 608806 480312 608812
rect 483216 605834 483244 619520
rect 483032 605806 483244 605834
rect 482652 580712 482704 580718
rect 482652 580654 482704 580660
rect 482744 580712 482796 580718
rect 482744 580654 482796 580660
rect 473728 567112 473780 567118
rect 473728 567054 473780 567060
rect 473912 567112 473964 567118
rect 473912 567054 473964 567060
rect 473740 365498 473768 567054
rect 473924 534750 473952 567054
rect 473912 534744 473964 534750
rect 473912 534686 473964 534692
rect 481824 500676 481876 500682
rect 481824 500618 481876 500624
rect 477776 485444 477828 485450
rect 477776 485386 477828 485392
rect 473728 365492 473780 365498
rect 473728 365434 473780 365440
rect 473636 365356 473688 365362
rect 473636 365298 473688 365304
rect 472624 191888 472676 191894
rect 472624 191830 472676 191836
rect 472636 111246 472664 191830
rect 473648 140486 473676 365298
rect 473636 140480 473688 140486
rect 473636 140422 473688 140428
rect 472624 111240 472676 111246
rect 472624 111182 472676 111188
rect 471888 107976 471940 107982
rect 471888 107918 471940 107924
rect 473740 78606 473768 365434
rect 477684 329316 477736 329322
rect 477684 329258 477736 329264
rect 475384 222420 475436 222426
rect 475384 222362 475436 222368
rect 473728 78600 473780 78606
rect 473728 78542 473780 78548
rect 475396 14074 475424 222362
rect 477696 126002 477724 329258
rect 477788 126138 477816 485386
rect 481732 329044 481784 329050
rect 481732 328986 481784 328992
rect 481744 314226 481772 328986
rect 481836 314362 481864 500618
rect 481824 314356 481876 314362
rect 481824 314298 481876 314304
rect 481732 314220 481784 314226
rect 481732 314162 481784 314168
rect 482664 130422 482692 580654
rect 482756 578950 482784 580654
rect 482744 578944 482796 578950
rect 482744 578886 482796 578892
rect 483032 325990 483060 605806
rect 484216 455456 484268 455462
rect 484216 455398 484268 455404
rect 483020 325984 483072 325990
rect 483020 325926 483072 325932
rect 483020 307828 483072 307834
rect 483020 307770 483072 307776
rect 483032 283354 483060 307770
rect 483756 301504 483808 301510
rect 483756 301446 483808 301452
rect 483020 283348 483072 283354
rect 483020 283290 483072 283296
rect 483768 257650 483796 301446
rect 483756 257644 483808 257650
rect 483756 257586 483808 257592
rect 483848 218816 483900 218822
rect 483848 218758 483900 218764
rect 483860 199986 483888 218758
rect 483848 199980 483900 199986
rect 483848 199922 483900 199928
rect 484228 157146 484256 455398
rect 485596 414112 485648 414118
rect 485596 414054 485648 414060
rect 485608 346866 485636 414054
rect 486976 364744 487028 364750
rect 486976 364686 487028 364692
rect 485412 346860 485464 346866
rect 485412 346802 485464 346808
rect 485596 346860 485648 346866
rect 485596 346802 485648 346808
rect 485424 217598 485452 346802
rect 486988 266830 487016 364686
rect 486976 266824 487028 266830
rect 486976 266766 487028 266772
rect 485596 266688 485648 266694
rect 485596 266630 485648 266636
rect 485608 256562 485636 266630
rect 485596 256556 485648 256562
rect 485596 256498 485648 256504
rect 485412 217592 485464 217598
rect 485412 217534 485464 217540
rect 484216 157140 484268 157146
rect 484216 157082 484268 157088
rect 486988 146946 487016 266766
rect 486976 146940 487028 146946
rect 486976 146882 487028 146888
rect 482652 130416 482704 130422
rect 482652 130358 482704 130364
rect 477776 126132 477828 126138
rect 477776 126074 477828 126080
rect 477684 125996 477736 126002
rect 477684 125938 477736 125944
rect 477696 120018 477724 125938
rect 477684 120012 477736 120018
rect 477684 119954 477736 119960
rect 489920 112192 489972 112198
rect 489920 112134 489972 112140
rect 480628 111648 480680 111654
rect 480628 111590 480680 111596
rect 480640 63510 480668 111590
rect 480628 63504 480680 63510
rect 480628 63446 480680 63452
rect 479432 37800 479484 37806
rect 479432 37742 479484 37748
rect 475384 14068 475436 14074
rect 475384 14010 475436 14016
rect 479444 13870 479472 37742
rect 489932 16574 489960 112134
rect 491312 108390 491340 619534
rect 492048 619426 492076 619534
rect 492190 619520 492302 620960
rect 495318 619520 495430 620960
rect 498262 619520 498374 620960
rect 492232 619426 492260 619520
rect 492048 619398 492260 619426
rect 495360 617574 495388 619520
rect 494060 617568 494112 617574
rect 494060 617510 494112 617516
rect 495348 617568 495400 617574
rect 495348 617510 495400 617516
rect 496174 617536 496230 617545
rect 492956 615528 493008 615534
rect 492956 615470 493008 615476
rect 492968 591258 492996 615470
rect 492956 591252 493008 591258
rect 492956 591194 493008 591200
rect 494072 111790 494100 617510
rect 496174 617471 496230 617480
rect 495438 613184 495494 613193
rect 495438 613119 495494 613128
rect 495452 612814 495480 613119
rect 495440 612808 495492 612814
rect 495440 612750 495492 612756
rect 495438 599584 495494 599593
rect 495438 599519 495494 599528
rect 495452 599010 495480 599519
rect 495440 599004 495492 599010
rect 495440 598946 495492 598952
rect 494336 591048 494388 591054
rect 494336 590990 494388 590996
rect 494348 469878 494376 590990
rect 495532 587308 495584 587314
rect 495532 587250 495584 587256
rect 495438 572928 495494 572937
rect 495438 572863 495494 572872
rect 495452 572762 495480 572863
rect 495440 572756 495492 572762
rect 495440 572698 495492 572704
rect 495438 554976 495494 554985
rect 495438 554911 495494 554920
rect 495452 554810 495480 554911
rect 495440 554804 495492 554810
rect 495440 554746 495492 554752
rect 495438 550352 495494 550361
rect 495438 550287 495494 550296
rect 495452 549302 495480 550287
rect 495440 549296 495492 549302
rect 495440 549238 495492 549244
rect 495438 546000 495494 546009
rect 495438 545935 495494 545944
rect 495452 545154 495480 545935
rect 495440 545148 495492 545154
rect 495440 545090 495492 545096
rect 495440 542360 495492 542366
rect 495440 542302 495492 542308
rect 495452 541385 495480 542302
rect 495438 541376 495494 541385
rect 495438 541311 495494 541320
rect 495438 537024 495494 537033
rect 495438 536959 495494 536968
rect 495452 536858 495480 536959
rect 495440 536852 495492 536858
rect 495440 536794 495492 536800
rect 495440 528556 495492 528562
rect 495440 528498 495492 528504
rect 495452 528057 495480 528498
rect 495438 528048 495494 528057
rect 495438 527983 495494 527992
rect 495438 510096 495494 510105
rect 495438 510031 495494 510040
rect 495452 509318 495480 510031
rect 495440 509312 495492 509318
rect 495440 509254 495492 509260
rect 495544 475726 495572 587250
rect 496082 532672 496138 532681
rect 496082 532607 496138 532616
rect 495532 475720 495584 475726
rect 495532 475662 495584 475668
rect 495624 475720 495676 475726
rect 495624 475662 495676 475668
rect 494336 469872 494388 469878
rect 494336 469814 494388 469820
rect 495438 469840 495494 469849
rect 495438 469775 495494 469784
rect 495452 469266 495480 469775
rect 495440 469260 495492 469266
rect 495440 469202 495492 469208
rect 495438 456512 495494 456521
rect 495438 456447 495494 456456
rect 495452 455462 495480 456447
rect 495440 455456 495492 455462
rect 495440 455398 495492 455404
rect 495438 442912 495494 442921
rect 495438 442847 495494 442856
rect 495452 441658 495480 442847
rect 495440 441652 495492 441658
rect 495440 441594 495492 441600
rect 495438 407280 495494 407289
rect 495438 407215 495494 407224
rect 495452 407182 495480 407215
rect 495440 407176 495492 407182
rect 495440 407118 495492 407124
rect 495440 402960 495492 402966
rect 495440 402902 495492 402908
rect 495452 402665 495480 402902
rect 495438 402656 495494 402665
rect 495438 402591 495494 402600
rect 495438 398304 495494 398313
rect 495438 398239 495494 398248
rect 495452 397594 495480 398239
rect 495440 397588 495492 397594
rect 495440 397530 495492 397536
rect 495440 385008 495492 385014
rect 495440 384950 495492 384956
rect 495452 384713 495480 384950
rect 495438 384704 495494 384713
rect 495438 384639 495494 384648
rect 495438 366752 495494 366761
rect 495438 366687 495494 366696
rect 495452 365770 495480 366687
rect 495440 365764 495492 365770
rect 495440 365706 495492 365712
rect 495438 362400 495494 362409
rect 495438 362335 495494 362344
rect 495452 361622 495480 362335
rect 495440 361616 495492 361622
rect 495440 361558 495492 361564
rect 495440 322924 495492 322930
rect 495440 322866 495492 322872
rect 495452 322153 495480 322866
rect 495438 322144 495494 322153
rect 495438 322079 495494 322088
rect 495440 313268 495492 313274
rect 495440 313210 495492 313216
rect 495452 313177 495480 313210
rect 495438 313168 495494 313177
rect 495438 313103 495494 313112
rect 495438 308544 495494 308553
rect 495438 308479 495494 308488
rect 495452 307834 495480 308479
rect 495440 307828 495492 307834
rect 495440 307770 495492 307776
rect 495636 304230 495664 475662
rect 495992 423700 496044 423706
rect 495992 423642 496044 423648
rect 496004 420617 496032 423642
rect 495990 420608 496046 420617
rect 495990 420543 496046 420552
rect 495624 304224 495676 304230
rect 495624 304166 495676 304172
rect 495440 300144 495492 300150
rect 495440 300086 495492 300092
rect 495452 299849 495480 300086
rect 495438 299840 495494 299849
rect 495438 299775 495494 299784
rect 495440 295316 495492 295322
rect 495440 295258 495492 295264
rect 495452 295225 495480 295258
rect 495438 295216 495494 295225
rect 495438 295151 495494 295160
rect 495440 286952 495492 286958
rect 495440 286894 495492 286900
rect 495452 286249 495480 286894
rect 495438 286240 495494 286249
rect 495438 286175 495494 286184
rect 495438 281888 495494 281897
rect 495438 281823 495494 281832
rect 495452 281586 495480 281823
rect 495440 281580 495492 281586
rect 495440 281522 495492 281528
rect 495990 272912 496046 272921
rect 495990 272847 496046 272856
rect 495438 268288 495494 268297
rect 495438 268223 495494 268232
rect 495452 267782 495480 268223
rect 495440 267776 495492 267782
rect 495440 267718 495492 267724
rect 495438 259312 495494 259321
rect 495438 259247 495494 259256
rect 495452 258126 495480 259247
rect 495440 258120 495492 258126
rect 495440 258062 495492 258068
rect 495440 251184 495492 251190
rect 495440 251126 495492 251132
rect 495452 250345 495480 251126
rect 495438 250336 495494 250345
rect 495438 250271 495494 250280
rect 496004 219638 496032 272847
rect 495992 219632 496044 219638
rect 495992 219574 496044 219580
rect 495438 219056 495494 219065
rect 495438 218991 495494 219000
rect 495452 218074 495480 218991
rect 495440 218068 495492 218074
rect 495440 218010 495492 218016
rect 495440 201476 495492 201482
rect 495440 201418 495492 201424
rect 495452 201113 495480 201418
rect 495438 201104 495494 201113
rect 495438 201039 495494 201048
rect 495440 197328 495492 197334
rect 495440 197270 495492 197276
rect 495452 196761 495480 197270
rect 495438 196752 495494 196761
rect 495438 196687 495494 196696
rect 495438 192128 495494 192137
rect 495438 192063 495494 192072
rect 495452 191894 495480 192063
rect 495440 191888 495492 191894
rect 495440 191830 495492 191836
rect 495438 187776 495494 187785
rect 495438 187711 495440 187720
rect 495492 187711 495494 187720
rect 495440 187682 495492 187688
rect 495440 175228 495492 175234
rect 495440 175170 495492 175176
rect 495452 174457 495480 175170
rect 495438 174448 495494 174457
rect 495438 174383 495494 174392
rect 495530 147520 495586 147529
rect 495530 147455 495586 147464
rect 495544 146946 495572 147455
rect 495532 146940 495584 146946
rect 495532 146882 495584 146888
rect 495440 143540 495492 143546
rect 495440 143482 495492 143488
rect 495452 142905 495480 143482
rect 495438 142896 495494 142905
rect 495438 142831 495494 142840
rect 495544 142154 495572 146882
rect 495452 142126 495572 142154
rect 495452 116618 495480 142126
rect 496096 118386 496124 532607
rect 496188 220697 496216 617471
rect 496358 604208 496414 604217
rect 496358 604143 496414 604152
rect 496266 595232 496322 595241
rect 496266 595167 496322 595176
rect 496280 295730 496308 595167
rect 496372 507958 496400 604143
rect 496360 507952 496412 507958
rect 496360 507894 496412 507900
rect 496360 507272 496412 507278
rect 496360 507214 496412 507220
rect 496372 478825 496400 507214
rect 496358 478816 496414 478825
rect 496358 478751 496414 478760
rect 496372 364614 496400 478751
rect 496450 474464 496506 474473
rect 496450 474399 496506 474408
rect 496360 364608 496412 364614
rect 496360 364550 496412 364556
rect 496358 358048 496414 358057
rect 496358 357983 496414 357992
rect 496268 295724 496320 295730
rect 496268 295666 496320 295672
rect 496266 277264 496322 277273
rect 496266 277199 496322 277208
rect 496280 240650 496308 277199
rect 496268 240644 496320 240650
rect 496268 240586 496320 240592
rect 496266 237008 496322 237017
rect 496266 236943 496322 236952
rect 496174 220688 496230 220697
rect 496174 220623 496230 220632
rect 496174 205728 496230 205737
rect 496174 205663 496230 205672
rect 496188 118590 496216 205663
rect 496280 118658 496308 236943
rect 496372 222902 496400 357983
rect 496360 222896 496412 222902
rect 496360 222838 496412 222844
rect 496360 217524 496412 217530
rect 496360 217466 496412 217472
rect 496372 183433 496400 217466
rect 496358 183424 496414 183433
rect 496358 183359 496414 183368
rect 496358 129568 496414 129577
rect 496358 129503 496414 129512
rect 496268 118652 496320 118658
rect 496268 118594 496320 118600
rect 496176 118584 496228 118590
rect 496176 118526 496228 118532
rect 496084 118380 496136 118386
rect 496084 118322 496136 118328
rect 495440 116612 495492 116618
rect 495440 116554 495492 116560
rect 494060 111784 494112 111790
rect 494060 111726 494112 111732
rect 495440 110832 495492 110838
rect 495440 110774 495492 110780
rect 491300 108384 491352 108390
rect 491300 108326 491352 108332
rect 493876 65544 493928 65550
rect 493876 65486 493928 65492
rect 489932 16546 490144 16574
rect 479432 13864 479484 13870
rect 479432 13806 479484 13812
rect 470048 4820 470100 4826
rect 470048 4762 470100 4768
rect 475476 3800 475528 3806
rect 475476 3742 475528 3748
rect 475488 480 475516 3742
rect 478418 3496 478474 3505
rect 478418 3431 478474 3440
rect 484492 3460 484544 3466
rect 478432 480 478460 3431
rect 484492 3402 484544 3408
rect 484504 480 484532 3402
rect 490116 490 490144 16546
rect 493888 3874 493916 65486
rect 495452 16574 495480 110774
rect 495530 102640 495586 102649
rect 495530 102575 495586 102584
rect 495544 102202 495572 102575
rect 495532 102196 495584 102202
rect 495532 102138 495584 102144
rect 495532 99272 495584 99278
rect 495532 99214 495584 99220
rect 495544 98297 495572 99214
rect 495530 98288 495586 98297
rect 495530 98223 495586 98232
rect 495532 93832 495584 93838
rect 495532 93774 495584 93780
rect 495544 93673 495572 93774
rect 495530 93664 495586 93673
rect 495530 93599 495586 93608
rect 495532 89684 495584 89690
rect 495532 89626 495584 89632
rect 495544 89321 495572 89626
rect 495530 89312 495586 89321
rect 495530 89247 495586 89256
rect 495532 63504 495584 63510
rect 495532 63446 495584 63452
rect 495544 62393 495572 63446
rect 495530 62384 495586 62393
rect 495530 62319 495586 62328
rect 496084 61124 496136 61130
rect 496084 61066 496136 61072
rect 495532 59220 495584 59226
rect 495532 59162 495584 59168
rect 495544 58041 495572 59162
rect 495530 58032 495586 58041
rect 495530 57967 495586 57976
rect 496096 55214 496124 61066
rect 496096 55186 496216 55214
rect 495532 45552 495584 45558
rect 495532 45494 495584 45500
rect 495544 44441 495572 45494
rect 495530 44432 495586 44441
rect 495530 44367 495586 44376
rect 496188 40089 496216 55186
rect 496372 43110 496400 129503
rect 496464 72282 496492 474399
rect 496542 451888 496598 451897
rect 496542 451823 496598 451832
rect 496556 432070 496584 451823
rect 496544 432064 496596 432070
rect 496544 432006 496596 432012
rect 496634 290864 496690 290873
rect 496634 290799 496690 290808
rect 496542 223680 496598 223689
rect 496542 223615 496598 223624
rect 496556 119270 496584 223615
rect 496648 223242 496676 290799
rect 496636 223236 496688 223242
rect 496636 223178 496688 223184
rect 496728 222352 496780 222358
rect 496728 222294 496780 222300
rect 496634 178800 496690 178809
rect 496634 178735 496690 178744
rect 496544 119264 496596 119270
rect 496544 119206 496596 119212
rect 496648 118522 496676 178735
rect 496740 169833 496768 222294
rect 496726 169824 496782 169833
rect 496726 169759 496782 169768
rect 496636 118516 496688 118522
rect 496636 118458 496688 118464
rect 496452 72276 496504 72282
rect 496452 72218 496504 72224
rect 496360 43104 496412 43110
rect 496360 43046 496412 43052
rect 496174 40080 496230 40089
rect 496174 40015 496230 40024
rect 495532 35896 495584 35902
rect 495532 35838 495584 35844
rect 495544 35465 495572 35838
rect 495530 35456 495586 35465
rect 495530 35391 495586 35400
rect 495532 23452 495584 23458
rect 495532 23394 495584 23400
rect 495544 22137 495572 23394
rect 495530 22128 495586 22137
rect 495530 22063 495586 22072
rect 495452 16546 496216 16574
rect 495440 13796 495492 13802
rect 495440 13738 495492 13744
rect 495452 13161 495480 13738
rect 495438 13152 495494 13161
rect 495438 13087 495494 13096
rect 495440 9580 495492 9586
rect 495440 9522 495492 9528
rect 495452 8809 495480 9522
rect 495438 8800 495494 8809
rect 495438 8735 495494 8744
rect 493876 3868 493928 3874
rect 493876 3810 493928 3816
rect 490392 598 490604 626
rect 490392 490 490420 598
rect 387678 -960 387790 480
rect 390622 -960 390734 480
rect 393566 -960 393678 480
rect 396694 -960 396806 480
rect 399638 -960 399750 480
rect 402766 -960 402878 480
rect 405710 -960 405822 480
rect 408838 -960 408950 480
rect 411782 -960 411894 480
rect 414910 -960 415022 480
rect 417854 -960 417966 480
rect 420982 -960 421094 480
rect 423926 -960 424038 480
rect 427054 -960 427166 480
rect 429998 -960 430110 480
rect 432942 -960 433054 480
rect 436070 -960 436182 480
rect 439014 -960 439126 480
rect 442142 -960 442254 480
rect 445086 -960 445198 480
rect 448214 -960 448326 480
rect 451158 -960 451270 480
rect 454286 -960 454398 480
rect 457230 -960 457342 480
rect 460358 -960 460470 480
rect 463302 -960 463414 480
rect 466430 -960 466542 480
rect 469374 -960 469486 480
rect 472318 -960 472430 480
rect 475446 -960 475558 480
rect 478390 -960 478502 480
rect 481518 -960 481630 480
rect 484462 -960 484574 480
rect 487590 -960 487702 480
rect 490116 462 490420 490
rect 490576 480 490604 598
rect 496188 490 496216 16546
rect 496360 15496 496412 15502
rect 496360 15438 496412 15444
rect 496372 9450 496400 15438
rect 496360 9444 496412 9450
rect 496360 9386 496412 9392
rect 499764 3256 499816 3262
rect 499764 3198 499816 3204
rect 496464 598 496676 626
rect 496464 490 496492 598
rect 490534 -960 490646 480
rect 493662 -960 493774 480
rect 496188 462 496492 490
rect 496648 480 496676 598
rect 499776 480 499804 3198
rect 496606 -960 496718 480
rect 499734 -960 499846 480
<< via2 >>
rect 3422 617752 3478 617808
rect 3054 608796 3110 608832
rect 3054 608776 3056 608796
rect 3056 608776 3108 608796
rect 3108 608776 3110 608796
rect 3422 604460 3424 604480
rect 3424 604460 3476 604480
rect 3476 604460 3478 604480
rect 3422 604424 3478 604460
rect 3514 599800 3570 599856
rect 2778 595448 2834 595504
rect 2778 586508 2780 586528
rect 2780 586508 2832 586528
rect 2832 586508 2834 586528
rect 2778 586472 2834 586508
rect 2778 577496 2834 577552
rect 2870 559544 2926 559600
rect 2778 555192 2834 555248
rect 3146 546216 3202 546272
rect 2870 541592 2926 541648
rect 3146 537240 3202 537296
rect 3330 514936 3386 514992
rect 3146 505960 3202 506016
rect 2778 497004 2834 497040
rect 2778 496984 2780 497004
rect 2780 496984 2832 497004
rect 2832 496984 2834 497004
rect 2778 479052 2834 479088
rect 2778 479032 2780 479052
rect 2780 479032 2832 479052
rect 2832 479032 2834 479052
rect 3330 461080 3386 461136
rect 3146 443128 3202 443184
rect 2962 402872 3018 402928
rect 2778 366968 2834 367024
rect 2870 205980 2872 206000
rect 2872 205980 2924 206000
rect 2924 205980 2926 206000
rect 2870 205944 2926 205980
rect 2778 120808 2834 120864
rect 3330 434152 3386 434208
rect 3238 429800 3294 429856
rect 3054 317736 3110 317792
rect 3330 425196 3386 425232
rect 3330 425176 3332 425196
rect 3332 425176 3384 425196
rect 3384 425176 3386 425196
rect 3330 407224 3386 407280
rect 3054 223896 3110 223952
rect 3330 246200 3386 246256
rect 3330 222536 3386 222592
rect 3238 201320 3294 201376
rect 3054 183404 3056 183424
rect 3056 183404 3108 183424
rect 3108 183404 3110 183424
rect 3054 183368 3110 183404
rect 3146 156712 3202 156768
rect 3146 117272 3202 117328
rect 2778 75928 2834 75984
rect 3146 66952 3202 67008
rect 2778 57976 2834 58032
rect 2778 53660 2780 53680
rect 2780 53660 2832 53680
rect 2832 53660 2834 53680
rect 2778 53624 2834 53660
rect 3330 187992 3386 188048
rect 3330 179016 3386 179072
rect 3330 161100 3332 161120
rect 3332 161100 3384 161120
rect 3384 161100 3386 161120
rect 3330 161064 3386 161100
rect 3330 138760 3386 138816
rect 3238 40296 3294 40352
rect 2778 8744 2834 8800
rect 3698 528264 3754 528320
rect 3882 519288 3938 519344
rect 3698 420824 3754 420880
rect 3606 389544 3662 389600
rect 3606 331336 3662 331392
rect 3606 322360 3662 322416
rect 3606 290808 3662 290864
rect 3606 273164 3608 273184
rect 3608 273164 3660 273184
rect 3660 273164 3662 273184
rect 3606 273128 3662 273164
rect 3606 268504 3662 268560
rect 3606 219272 3662 219328
rect 3606 214920 3662 214976
rect 3790 416200 3846 416256
rect 3790 384920 3846 384976
rect 3698 117952 3754 118008
rect 3882 264152 3938 264208
rect 3882 255176 3938 255232
rect 3790 84904 3846 84960
rect 3514 80552 3570 80608
rect 3422 35672 3478 35728
rect 3422 17720 3478 17776
rect 3330 8608 3386 8664
rect 4158 308760 4214 308816
rect 4066 152088 4122 152144
rect 3974 143112 4030 143168
rect 4066 134136 4122 134192
rect 4066 129784 4122 129840
rect 3974 125160 4030 125216
rect 4066 111832 4122 111888
rect 4066 44648 4122 44704
rect 5446 220088 5502 220144
rect 3422 7928 3478 7984
rect 5814 118224 5870 118280
rect 7010 158752 7066 158808
rect 6918 149096 6974 149152
rect 7378 197784 7434 197840
rect 7470 178880 7526 178936
rect 7378 168408 7434 168464
rect 7286 113872 7342 113928
rect 7562 149096 7618 149152
rect 7470 68856 7526 68912
rect 7378 59200 7434 59256
rect 7194 49544 7250 49600
rect 7654 139712 7710 139768
rect 7562 39888 7618 39944
rect 7654 30232 7710 30288
rect 8022 208256 8078 208312
rect 7930 108568 7986 108624
rect 8022 98776 8078 98832
rect 8022 88984 8078 89040
rect 8206 188944 8262 189000
rect 8206 129920 8262 129976
rect 8114 78512 8170 78568
rect 8114 59200 8170 59256
rect 8206 20440 8262 20496
rect 8942 121352 8998 121408
rect 9126 109112 9182 109168
rect 9494 217776 9550 217832
rect 9126 9424 9182 9480
rect 32310 493060 32366 493096
rect 32310 493040 32312 493060
rect 32312 493040 32364 493060
rect 32364 493040 32366 493060
rect 32402 492632 32458 492688
rect 50158 599020 50160 599040
rect 50160 599020 50212 599040
rect 50212 599020 50214 599040
rect 50158 598984 50214 599020
rect 39394 381012 39396 381032
rect 39396 381012 39448 381032
rect 39448 381012 39450 381032
rect 39394 380976 39450 381012
rect 38842 333260 38898 333296
rect 38842 333240 38844 333260
rect 38844 333240 38896 333260
rect 38896 333240 38898 333260
rect 47674 435004 47676 435024
rect 47676 435004 47728 435024
rect 47728 435004 47730 435024
rect 47674 434968 47730 435004
rect 48042 434696 48098 434752
rect 34794 219952 34850 220008
rect 42062 219952 42118 220008
rect 49974 219952 50030 220008
rect 55310 409964 55366 410000
rect 75918 566072 75974 566128
rect 55310 409944 55312 409964
rect 55312 409944 55364 409964
rect 55364 409944 55366 409964
rect 55034 220516 55090 220552
rect 55034 220496 55036 220516
rect 55036 220496 55088 220516
rect 55088 220496 55090 220516
rect 54666 219952 54722 220008
rect 76286 565800 76342 565856
rect 67362 400596 67364 400616
rect 67364 400596 67416 400616
rect 67416 400596 67418 400616
rect 67362 400560 67418 400596
rect 67546 400560 67602 400616
rect 67638 400288 67694 400344
rect 62486 236172 62488 236192
rect 62488 236172 62540 236192
rect 62540 236172 62542 236192
rect 62486 236136 62542 236172
rect 61474 236000 61530 236056
rect 61842 222264 61898 222320
rect 68282 219952 68338 220008
rect 75182 222264 75238 222320
rect 77758 219680 77814 219736
rect 92386 616800 92442 616856
rect 93766 473492 93768 473512
rect 93768 473492 93820 473512
rect 93820 473492 93822 473512
rect 93766 473456 93822 473492
rect 91466 433336 91522 433392
rect 88798 383968 88854 384024
rect 90638 356496 90694 356552
rect 92938 288108 92994 288144
rect 92938 288088 92940 288108
rect 92940 288088 92992 288108
rect 92992 288088 92994 288108
rect 93122 288108 93178 288144
rect 93122 288088 93124 288108
rect 93124 288088 93176 288108
rect 93176 288088 93178 288108
rect 79322 220632 79378 220688
rect 79414 219952 79470 220008
rect 94502 219952 94558 220008
rect 98734 263608 98790 263664
rect 100942 224440 100998 224496
rect 101402 219952 101458 220008
rect 87786 219408 87842 219464
rect 96618 219408 96674 219464
rect 112350 446956 112406 446992
rect 112350 446936 112352 446956
rect 112352 446936 112404 446956
rect 112404 446936 112406 446956
rect 103518 384140 103520 384160
rect 103520 384140 103572 384160
rect 103572 384140 103574 384160
rect 103518 384104 103574 384140
rect 112166 295568 112222 295624
rect 103426 266872 103482 266928
rect 103426 248376 103482 248432
rect 103426 238584 103482 238640
rect 103426 229064 103482 229120
rect 103426 228928 103482 228984
rect 103426 224848 103482 224904
rect 112810 410488 112866 410544
rect 119986 541476 120042 541512
rect 119986 541456 119988 541476
rect 119988 541456 120040 541476
rect 120040 541456 120042 541476
rect 119618 414024 119674 414080
rect 114466 295568 114522 295624
rect 123298 541628 123300 541648
rect 123300 541628 123352 541648
rect 123352 541628 123354 541648
rect 123298 541592 123354 541628
rect 132590 384276 132592 384296
rect 132592 384276 132644 384296
rect 132644 384276 132646 384296
rect 132590 384240 132646 384276
rect 125322 261160 125378 261216
rect 125874 260908 125930 260944
rect 125874 260888 125876 260908
rect 125876 260888 125928 260908
rect 125928 260888 125930 260908
rect 123390 220632 123446 220688
rect 114926 219408 114982 219464
rect 130474 261160 130530 261216
rect 131578 260908 131634 260944
rect 131578 260888 131580 260908
rect 131580 260888 131632 260908
rect 131632 260888 131634 260908
rect 140778 307012 140834 307048
rect 140778 306992 140780 307012
rect 140780 306992 140832 307012
rect 140832 306992 140834 307012
rect 135626 227024 135682 227080
rect 136546 227060 136548 227080
rect 136548 227060 136600 227080
rect 136600 227060 136602 227080
rect 136546 227024 136602 227060
rect 137190 226616 137246 226672
rect 152370 442992 152426 443048
rect 143078 365372 143080 365392
rect 143080 365372 143132 365392
rect 143132 365372 143134 365392
rect 143078 365336 143134 365372
rect 134522 219952 134578 220008
rect 177210 616256 177266 616312
rect 157430 543788 157486 543824
rect 157430 543768 157432 543788
rect 157432 543768 157484 543788
rect 157484 543768 157486 543788
rect 159086 539552 159142 539608
rect 153474 229780 153476 229800
rect 153476 229780 153528 229800
rect 153528 229780 153530 229800
rect 153474 229744 153530 229780
rect 159270 273808 159326 273864
rect 159086 220224 159142 220280
rect 154026 219952 154082 220008
rect 167458 228268 167514 228304
rect 167458 228248 167460 228268
rect 167460 228248 167512 228268
rect 167512 228248 167514 228268
rect 167366 228148 167368 228168
rect 167368 228148 167420 228168
rect 167420 228148 167422 228168
rect 167366 228112 167422 228148
rect 177210 383852 177266 383888
rect 177210 383832 177212 383852
rect 177212 383832 177264 383852
rect 177264 383832 177266 383852
rect 175830 228148 175832 228168
rect 175832 228148 175884 228168
rect 175884 228148 175886 228168
rect 175830 228112 175886 228148
rect 180062 362500 180118 362536
rect 180062 362480 180064 362500
rect 180064 362480 180116 362500
rect 180116 362480 180118 362500
rect 190366 499568 190422 499624
rect 205454 596400 205510 596456
rect 205914 596300 205916 596320
rect 205916 596300 205968 596320
rect 205968 596300 205970 596320
rect 201498 583752 201554 583808
rect 198278 470600 198334 470656
rect 194598 353404 194600 353424
rect 194600 353404 194652 353424
rect 194652 353404 194654 353424
rect 194598 353368 194654 353404
rect 180890 259140 180946 259176
rect 180890 259120 180892 259140
rect 180892 259120 180944 259140
rect 180944 259120 180946 259140
rect 180798 258576 180854 258632
rect 162766 219544 162822 219600
rect 161294 219408 161350 219464
rect 187146 219952 187202 220008
rect 193770 219952 193826 220008
rect 205914 596264 205970 596300
rect 208582 498092 208638 498128
rect 208582 498072 208584 498092
rect 208584 498072 208636 498092
rect 208636 498072 208638 498092
rect 207386 262420 207388 262440
rect 207388 262420 207440 262440
rect 207440 262420 207442 262440
rect 207386 262384 207442 262420
rect 214746 369824 214802 369880
rect 231858 616800 231914 616856
rect 234802 616800 234858 616856
rect 240874 616800 240930 616856
rect 228454 606056 228510 606112
rect 218702 337592 218758 337648
rect 214378 222400 214434 222456
rect 207386 222264 207442 222320
rect 209042 220788 209098 220824
rect 209042 220768 209044 220788
rect 209044 220768 209096 220788
rect 209096 220768 209098 220788
rect 213182 220396 213184 220416
rect 213184 220396 213236 220416
rect 213236 220396 213238 220416
rect 213182 220360 213238 220396
rect 205178 219580 205180 219600
rect 205180 219580 205232 219600
rect 205232 219580 205234 219600
rect 205178 219544 205234 219580
rect 167918 219408 167974 219464
rect 173990 219408 174046 219464
rect 181166 219408 181222 219464
rect 219806 254788 219862 254824
rect 219806 254768 219808 254788
rect 219808 254768 219860 254788
rect 219860 254768 219862 254788
rect 219254 254668 219256 254688
rect 219256 254668 219308 254688
rect 219308 254668 219310 254688
rect 219254 254632 219310 254668
rect 231030 337320 231086 337376
rect 229098 267824 229154 267880
rect 259090 615576 259146 615632
rect 233698 371728 233754 371784
rect 226982 219952 227038 220008
rect 240322 232484 240378 232520
rect 240322 232464 240324 232484
rect 240324 232464 240376 232484
rect 240376 232464 240378 232484
rect 240138 222536 240194 222592
rect 235262 219952 235318 220008
rect 240138 219680 240194 219736
rect 234158 219408 234214 219464
rect 220266 219272 220322 219328
rect 248234 273808 248290 273864
rect 262770 525292 262826 525328
rect 262770 525272 262772 525292
rect 262772 525272 262824 525292
rect 262824 525272 262826 525292
rect 262678 525172 262680 525192
rect 262680 525172 262732 525192
rect 262732 525172 262734 525192
rect 255962 223236 256018 223272
rect 255962 223216 255964 223236
rect 255964 223216 256016 223236
rect 256016 223216 256018 223236
rect 262678 525136 262734 525172
rect 263690 436056 263746 436112
rect 259182 220652 259238 220688
rect 261114 300872 261170 300928
rect 260746 223236 260802 223272
rect 260746 223216 260748 223236
rect 260748 223216 260800 223236
rect 260800 223216 260802 223236
rect 259182 220632 259184 220652
rect 259184 220632 259236 220652
rect 259236 220632 259238 220652
rect 253386 219952 253442 220008
rect 257710 219816 257766 219872
rect 274178 616120 274234 616176
rect 268290 553424 268346 553480
rect 268566 553424 268622 553480
rect 281630 432132 281686 432168
rect 281630 432112 281632 432132
rect 281632 432112 281684 432132
rect 281684 432112 281686 432132
rect 282734 432012 282736 432032
rect 282736 432012 282788 432032
rect 282788 432012 282790 432032
rect 282734 431976 282790 432012
rect 274454 380452 274510 380488
rect 274454 380432 274456 380452
rect 274456 380432 274508 380452
rect 274508 380432 274510 380452
rect 282274 324980 282276 325000
rect 282276 324980 282328 325000
rect 282328 324980 282330 325000
rect 282274 324944 282330 324980
rect 273626 287020 273682 287056
rect 273626 287000 273628 287020
rect 273628 287000 273680 287020
rect 273680 287000 273682 287020
rect 273994 285640 274050 285696
rect 283378 610000 283434 610056
rect 295338 616800 295394 616856
rect 289818 518644 289820 518664
rect 289820 518644 289872 518664
rect 289872 518644 289874 518664
rect 289818 518608 289874 518644
rect 291106 518764 291162 518800
rect 291106 518744 291108 518764
rect 291108 518744 291160 518764
rect 291160 518744 291162 518764
rect 264978 219836 265034 219872
rect 303158 249872 303214 249928
rect 289634 223624 289690 223680
rect 280526 219952 280582 220008
rect 264978 219816 264980 219836
rect 264980 219816 265032 219836
rect 265032 219816 265034 219836
rect 266634 219816 266690 219872
rect 273258 219408 273314 219464
rect 293222 219408 293278 219464
rect 244922 219272 244978 219328
rect 9862 111968 9918 112024
rect 43534 120672 43590 120728
rect 96434 120672 96490 120728
rect 103150 120672 103206 120728
rect 116398 120672 116454 120728
rect 34978 119992 35034 120048
rect 35162 119856 35218 119912
rect 35346 119468 35402 119504
rect 35346 119448 35348 119468
rect 35348 119448 35400 119468
rect 35400 119448 35402 119468
rect 34886 119312 34942 119368
rect 34610 119060 34666 119096
rect 34610 119040 34612 119060
rect 34612 119040 34664 119060
rect 34664 119040 34666 119060
rect 34794 118904 34850 118960
rect 34886 118804 34888 118824
rect 34888 118804 34940 118824
rect 34940 118804 34942 118824
rect 34886 118768 34942 118804
rect 29734 117816 29790 117872
rect 32494 113892 32550 113928
rect 32494 113872 32496 113892
rect 32496 113872 32548 113892
rect 32548 113872 32550 113892
rect 35070 111968 35126 112024
rect 38750 119992 38806 120048
rect 48134 119176 48190 119232
rect 38842 119040 38898 119096
rect 49882 118496 49938 118552
rect 56230 118088 56286 118144
rect 63498 119992 63554 120048
rect 63682 119992 63738 120048
rect 64050 119312 64106 119368
rect 76378 118088 76434 118144
rect 36634 117408 36690 117464
rect 49882 117408 49938 117464
rect 62762 117408 62818 117464
rect 83002 117408 83058 117464
rect 109130 118360 109186 118416
rect 122194 117816 122250 117872
rect 145654 119040 145710 119096
rect 145746 118768 145802 118824
rect 142342 118088 142398 118144
rect 161018 119992 161074 120048
rect 157522 119040 157578 119096
rect 162490 119856 162546 119912
rect 135994 117408 136050 117464
rect 149518 117408 149574 117464
rect 155590 117408 155646 117464
rect 162214 117408 162270 117464
rect 69386 114416 69442 114472
rect 41694 111968 41750 112024
rect 61566 112104 61622 112160
rect 68190 112104 68246 112160
rect 54942 111968 54998 112024
rect 74814 111968 74870 112024
rect 88062 111968 88118 112024
rect 94686 111968 94742 112024
rect 101310 111968 101366 112024
rect 96894 110608 96950 110664
rect 160926 112784 160982 112840
rect 107934 112512 107990 112568
rect 115110 112104 115166 112160
rect 141054 112512 141110 112568
rect 134430 112104 134486 112160
rect 132774 111580 132830 111616
rect 132774 111560 132776 111580
rect 132776 111560 132828 111580
rect 132828 111560 132830 111580
rect 135718 110880 135774 110936
rect 137190 110508 137192 110528
rect 137192 110508 137244 110528
rect 137244 110508 137246 110528
rect 137190 110472 137246 110508
rect 147678 112104 147734 112160
rect 154302 112104 154358 112160
rect 167550 112784 167606 112840
rect 172702 119992 172758 120048
rect 168746 118224 168802 118280
rect 175922 117408 175978 117464
rect 174174 111832 174230 111888
rect 170218 111152 170274 111208
rect 168378 110764 168434 110800
rect 168378 110744 168380 110764
rect 168380 110744 168432 110764
rect 168432 110744 168434 110764
rect 168102 110472 168158 110528
rect 180798 112240 180854 112296
rect 180614 111696 180670 111752
rect 179510 111424 179566 111480
rect 179326 111288 179382 111344
rect 188986 118224 189042 118280
rect 215758 119720 215814 119776
rect 215574 119584 215630 119640
rect 216034 119448 216090 119504
rect 215850 119040 215906 119096
rect 216586 119040 216642 119096
rect 209134 118124 209136 118144
rect 209136 118124 209188 118144
rect 209188 118124 209190 118144
rect 209134 118088 209190 118124
rect 182638 117408 182694 117464
rect 188986 117408 189042 117464
rect 195334 117408 195390 117464
rect 202234 117408 202290 117464
rect 209870 115776 209926 115832
rect 187422 113056 187478 113112
rect 194046 113056 194102 113112
rect 181258 111560 181314 111616
rect 182638 111288 182694 111344
rect 183466 111288 183522 111344
rect 181810 111172 181866 111208
rect 181810 111152 181812 111172
rect 181812 111152 181864 111172
rect 181864 111152 181866 111172
rect 183190 111152 183246 111208
rect 182638 110472 182694 110528
rect 190458 110508 190460 110528
rect 190460 110508 190512 110528
rect 190512 110508 190514 110528
rect 190458 110472 190514 110508
rect 200670 112648 200726 112704
rect 194414 111016 194470 111072
rect 207294 111832 207350 111888
rect 220542 113056 220598 113112
rect 213918 112648 213974 112704
rect 213642 111424 213698 111480
rect 214470 111288 214526 111344
rect 214654 111016 214710 111072
rect 214562 110880 214618 110936
rect 214746 110880 214802 110936
rect 238758 119176 238814 119232
rect 235630 118496 235686 118552
rect 241702 118224 241758 118280
rect 253938 119620 253940 119640
rect 253940 119620 253992 119640
rect 253992 119620 253994 119640
rect 253938 119584 253994 119620
rect 254490 119620 254492 119640
rect 254492 119620 254544 119640
rect 254544 119620 254546 119640
rect 254490 119584 254546 119620
rect 254214 119312 254270 119368
rect 261482 118632 261538 118688
rect 254858 118360 254914 118416
rect 268474 118088 268530 118144
rect 248878 117952 248934 118008
rect 228822 117408 228878 117464
rect 235630 117408 235686 117464
rect 241702 117408 241758 117464
rect 227166 113056 227222 113112
rect 273258 113056 273314 113112
rect 222382 111152 222438 111208
rect 222198 110472 222254 110528
rect 247038 112376 247094 112432
rect 233790 111968 233846 112024
rect 231858 111172 231914 111208
rect 231858 111152 231860 111172
rect 231860 111152 231912 111172
rect 231912 111152 231914 111172
rect 240414 111832 240470 111888
rect 253662 111832 253718 111888
rect 273166 110608 273222 110664
rect 281998 117408 282054 117464
rect 290462 119856 290518 119912
rect 289726 119468 289782 119504
rect 289726 119448 289728 119468
rect 289728 119448 289780 119468
rect 289780 119448 289782 119468
rect 292118 119448 292174 119504
rect 295154 117716 295156 117736
rect 295156 117716 295208 117736
rect 295208 117716 295210 117736
rect 295154 117680 295210 117716
rect 287978 117272 288034 117328
rect 286782 112512 286838 112568
rect 280158 111832 280214 111888
rect 273810 110744 273866 110800
rect 273626 110472 273682 110528
rect 293406 111832 293462 111888
rect 88154 109384 88210 109440
rect 29642 10648 29698 10704
rect 49882 10648 49938 10704
rect 56138 10648 56194 10704
rect 62762 10648 62818 10704
rect 36542 9832 36598 9888
rect 35530 9324 35532 9344
rect 35532 9324 35584 9344
rect 35584 9324 35586 9344
rect 35530 9288 35586 9324
rect 43166 8064 43222 8120
rect 11978 3304 12034 3360
rect 36266 3440 36322 3496
rect 122378 10648 122434 10704
rect 155498 10648 155554 10704
rect 162122 10648 162178 10704
rect 175922 10648 175978 10704
rect 65154 9444 65210 9480
rect 65154 9424 65156 9444
rect 65156 9424 65208 9444
rect 65208 9424 65210 9444
rect 66166 9424 66222 9480
rect 66166 9152 66222 9208
rect 51354 3440 51410 3496
rect 82910 9832 82966 9888
rect 77298 9596 77300 9616
rect 77300 9596 77352 9616
rect 77352 9596 77354 9616
rect 77298 9560 77354 9596
rect 77850 9580 77906 9616
rect 77850 9560 77852 9580
rect 77852 9560 77904 9580
rect 77904 9560 77906 9580
rect 78586 9596 78588 9616
rect 78588 9596 78640 9616
rect 78640 9596 78642 9616
rect 78586 9560 78642 9596
rect 79046 9424 79102 9480
rect 79230 9460 79232 9480
rect 79232 9460 79284 9480
rect 79284 9460 79286 9480
rect 79230 9424 79286 9460
rect 77942 9324 77944 9344
rect 77944 9324 77996 9344
rect 77996 9324 77998 9344
rect 77942 9288 77998 9324
rect 78862 9288 78918 9344
rect 77114 8880 77170 8936
rect 76286 8200 76342 8256
rect 88430 8880 88486 8936
rect 88614 8744 88670 8800
rect 88338 8472 88394 8528
rect 82910 7928 82966 7984
rect 95146 9580 95202 9616
rect 95146 9560 95148 9580
rect 95148 9560 95200 9580
rect 95200 9560 95202 9580
rect 96158 7928 96214 7984
rect 72698 3440 72754 3496
rect 109406 8064 109462 8120
rect 116490 9580 116546 9616
rect 116490 9560 116492 9580
rect 116492 9560 116544 9580
rect 116544 9560 116546 9580
rect 116030 7928 116086 7984
rect 102782 7792 102838 7848
rect 102874 3984 102930 4040
rect 100114 3712 100170 3768
rect 99930 3440 99986 3496
rect 100114 3440 100170 3496
rect 106002 3712 106058 3768
rect 135902 9832 135958 9888
rect 142250 9832 142306 9888
rect 148046 9016 148102 9072
rect 149518 10104 149574 10160
rect 168470 9696 168526 9752
rect 152554 8880 152610 8936
rect 168930 9716 168986 9752
rect 168930 9696 168932 9716
rect 168932 9696 168984 9716
rect 168984 9696 168986 9716
rect 168746 9580 168802 9616
rect 168746 9560 168748 9580
rect 168748 9560 168800 9580
rect 168800 9560 168802 9580
rect 169298 9580 169354 9616
rect 169298 9560 169300 9580
rect 169300 9560 169352 9580
rect 169352 9560 169354 9580
rect 169022 8064 169078 8120
rect 182638 10648 182694 10704
rect 188986 10648 189042 10704
rect 195242 10648 195298 10704
rect 202234 10648 202290 10704
rect 208858 10648 208914 10704
rect 228362 10648 228418 10704
rect 235630 10648 235686 10704
rect 185766 9560 185822 9616
rect 244554 10240 244610 10296
rect 241702 10104 241758 10160
rect 240046 9152 240102 9208
rect 239862 9016 239918 9072
rect 239862 8608 239918 8664
rect 244278 8744 244334 8800
rect 248142 9424 248198 9480
rect 248878 10648 248934 10704
rect 254858 10648 254914 10704
rect 261482 10648 261538 10704
rect 268750 10648 268806 10704
rect 274730 10648 274786 10704
rect 281998 10648 282054 10704
rect 287978 10648 288034 10704
rect 294602 10648 294658 10704
rect 272062 9560 272118 9616
rect 270866 9288 270922 9344
rect 270682 9152 270738 9208
rect 270958 8880 271014 8936
rect 272154 9016 272210 9072
rect 273166 9580 273222 9616
rect 273166 9560 273168 9580
rect 273168 9560 273220 9580
rect 273220 9560 273222 9580
rect 277766 9560 277822 9616
rect 273442 9424 273498 9480
rect 273810 9288 273866 9344
rect 277582 8880 277638 8936
rect 278134 9016 278190 9072
rect 272338 8336 272394 8392
rect 124034 3712 124090 3768
rect 142250 3032 142306 3088
rect 178682 3984 178738 4040
rect 151450 3848 151506 3904
rect 175554 3576 175610 3632
rect 169482 3168 169538 3224
rect 211986 3712 212042 3768
rect 221002 3440 221058 3496
rect 242162 3576 242218 3632
rect 263506 3984 263562 4040
rect 251362 3440 251418 3496
rect 266450 3712 266506 3768
rect 281538 3576 281594 3632
rect 310610 45872 310666 45928
rect 311714 220088 311770 220144
rect 312082 205128 312138 205184
rect 312174 185544 312230 185600
rect 312082 165960 312138 166016
rect 311990 85484 311992 85504
rect 311992 85484 312044 85504
rect 312044 85484 312046 85504
rect 311990 85448 312046 85484
rect 311898 17856 311954 17912
rect 311898 16904 311954 16960
rect 312174 156168 312230 156224
rect 312450 214920 312506 214976
rect 312634 214920 312690 214976
rect 312542 205128 312598 205184
rect 312450 185544 312506 185600
rect 312358 175752 312414 175808
rect 312266 146376 312322 146432
rect 312266 126792 312322 126848
rect 312082 55936 312138 55992
rect 312910 195336 312966 195392
rect 312726 146376 312782 146432
rect 312818 136584 312874 136640
rect 312634 105576 312690 105632
rect 312542 95104 312598 95160
rect 312450 75792 312506 75848
rect 312358 66136 312414 66192
rect 312450 55936 312506 55992
rect 312726 36660 312728 36680
rect 312728 36660 312780 36680
rect 312780 36660 312782 36680
rect 312726 36624 312782 36660
rect 312542 27240 312598 27296
rect 312266 17856 312322 17912
rect 313922 3440 313978 3496
rect 318246 220224 318302 220280
rect 373998 220496 374054 220552
rect 375378 3576 375434 3632
rect 415490 3304 415546 3360
rect 496174 617480 496230 617536
rect 495438 613128 495494 613184
rect 495438 599528 495494 599584
rect 495438 572872 495494 572928
rect 495438 554920 495494 554976
rect 495438 550296 495494 550352
rect 495438 545944 495494 546000
rect 495438 541320 495494 541376
rect 495438 536968 495494 537024
rect 495438 527992 495494 528048
rect 495438 510040 495494 510096
rect 496082 532616 496138 532672
rect 495438 469784 495494 469840
rect 495438 456456 495494 456512
rect 495438 442856 495494 442912
rect 495438 407224 495494 407280
rect 495438 402600 495494 402656
rect 495438 398248 495494 398304
rect 495438 384648 495494 384704
rect 495438 366696 495494 366752
rect 495438 362344 495494 362400
rect 495438 322088 495494 322144
rect 495438 313112 495494 313168
rect 495438 308488 495494 308544
rect 495990 420552 496046 420608
rect 495438 299784 495494 299840
rect 495438 295160 495494 295216
rect 495438 286184 495494 286240
rect 495438 281832 495494 281888
rect 495990 272856 496046 272912
rect 495438 268232 495494 268288
rect 495438 259256 495494 259312
rect 495438 250280 495494 250336
rect 495438 219000 495494 219056
rect 495438 201048 495494 201104
rect 495438 196696 495494 196752
rect 495438 192072 495494 192128
rect 495438 187740 495494 187776
rect 495438 187720 495440 187740
rect 495440 187720 495492 187740
rect 495492 187720 495494 187740
rect 495438 174392 495494 174448
rect 495530 147464 495586 147520
rect 495438 142840 495494 142896
rect 496358 604152 496414 604208
rect 496266 595176 496322 595232
rect 496358 478760 496414 478816
rect 496450 474408 496506 474464
rect 496358 357992 496414 358048
rect 496266 277208 496322 277264
rect 496266 236952 496322 237008
rect 496174 220632 496230 220688
rect 496174 205672 496230 205728
rect 496358 183368 496414 183424
rect 496358 129512 496414 129568
rect 478418 3440 478474 3496
rect 495530 102584 495586 102640
rect 495530 98232 495586 98288
rect 495530 93608 495586 93664
rect 495530 89256 495586 89312
rect 495530 62328 495586 62384
rect 495530 57976 495586 58032
rect 495530 44376 495586 44432
rect 496542 451832 496598 451888
rect 496634 290808 496690 290864
rect 496542 223624 496598 223680
rect 496634 178744 496690 178800
rect 496726 169768 496782 169824
rect 496174 40024 496230 40080
rect 495530 35400 495586 35456
rect 495530 22072 495586 22128
rect 495438 13096 495494 13152
rect 495438 8744 495494 8800
<< metal3 >>
rect -960 617810 480 617900
rect 3417 617810 3483 617813
rect -960 617808 3483 617810
rect -960 617752 3422 617808
rect 3478 617752 3483 617808
rect -960 617750 3483 617752
rect -960 617660 480 617750
rect 3417 617747 3483 617750
rect 496169 617538 496235 617541
rect 499520 617538 500960 617628
rect 496169 617536 500960 617538
rect 496169 617480 496174 617536
rect 496230 617480 500960 617536
rect 496169 617478 500960 617480
rect 496169 617475 496235 617478
rect 499520 617388 500960 617478
rect 90766 616796 90772 616860
rect 90836 616858 90842 616860
rect 92381 616858 92447 616861
rect 90836 616856 92447 616858
rect 90836 616800 92386 616856
rect 92442 616800 92447 616856
rect 90836 616798 92447 616800
rect 90836 616796 90842 616798
rect 92381 616795 92447 616798
rect 231853 616858 231919 616861
rect 232446 616858 232452 616860
rect 231853 616856 232452 616858
rect 231853 616800 231858 616856
rect 231914 616800 232452 616856
rect 231853 616798 232452 616800
rect 231853 616795 231919 616798
rect 232446 616796 232452 616798
rect 232516 616796 232522 616860
rect 234654 616796 234660 616860
rect 234724 616858 234730 616860
rect 234797 616858 234863 616861
rect 234724 616856 234863 616858
rect 234724 616800 234802 616856
rect 234858 616800 234863 616856
rect 234724 616798 234863 616800
rect 234724 616796 234730 616798
rect 234797 616795 234863 616798
rect 240869 616858 240935 616861
rect 295333 616860 295399 616861
rect 246246 616858 246252 616860
rect 240869 616856 246252 616858
rect 240869 616800 240874 616856
rect 240930 616800 246252 616856
rect 240869 616798 246252 616800
rect 240869 616795 240935 616798
rect 246246 616796 246252 616798
rect 246316 616796 246322 616860
rect 295333 616856 295380 616860
rect 295444 616858 295450 616860
rect 295333 616800 295338 616856
rect 295333 616796 295380 616800
rect 295444 616798 295490 616858
rect 295444 616796 295450 616798
rect 295333 616795 295399 616796
rect 177205 616314 177271 616317
rect 184054 616314 184060 616316
rect 177205 616312 184060 616314
rect 177205 616256 177210 616312
rect 177266 616256 184060 616312
rect 177205 616254 184060 616256
rect 177205 616251 177271 616254
rect 184054 616252 184060 616254
rect 184124 616252 184130 616316
rect 105486 616116 105492 616180
rect 105556 616178 105562 616180
rect 274173 616178 274239 616181
rect 105556 616176 274239 616178
rect 105556 616120 274178 616176
rect 274234 616120 274239 616176
rect 105556 616118 274239 616120
rect 105556 616116 105562 616118
rect 274173 616115 274239 616118
rect 258022 615572 258028 615636
rect 258092 615634 258098 615636
rect 259085 615634 259151 615637
rect 258092 615632 259151 615634
rect 258092 615576 259090 615632
rect 259146 615576 259151 615632
rect 258092 615574 259151 615576
rect 258092 615572 258098 615574
rect 259085 615571 259151 615574
rect -960 613308 480 613548
rect 495433 613186 495499 613189
rect 499520 613186 500960 613276
rect 495433 613184 500960 613186
rect 495433 613128 495438 613184
rect 495494 613128 500960 613184
rect 495433 613126 500960 613128
rect 495433 613123 495499 613126
rect 499520 613036 500960 613126
rect 283373 610060 283439 610061
rect 283373 610056 283420 610060
rect 283484 610058 283490 610060
rect 283373 610000 283378 610056
rect 283373 609996 283420 610000
rect 283484 609998 283530 610058
rect 283484 609996 283490 609998
rect 283373 609995 283439 609996
rect -960 608834 480 608924
rect 3049 608834 3115 608837
rect -960 608832 3115 608834
rect -960 608776 3054 608832
rect 3110 608776 3115 608832
rect -960 608774 3115 608776
rect -960 608684 480 608774
rect 3049 608771 3115 608774
rect 499520 608412 500960 608652
rect 228449 606114 228515 606117
rect 228582 606114 228588 606116
rect 228449 606112 228588 606114
rect 228449 606056 228454 606112
rect 228510 606056 228588 606112
rect 228449 606054 228588 606056
rect 228449 606051 228515 606054
rect 228582 606052 228588 606054
rect 228652 606052 228658 606116
rect -960 604482 480 604572
rect 3417 604482 3483 604485
rect -960 604480 3483 604482
rect -960 604424 3422 604480
rect 3478 604424 3483 604480
rect -960 604422 3483 604424
rect -960 604332 480 604422
rect 3417 604419 3483 604422
rect 496353 604210 496419 604213
rect 499520 604210 500960 604300
rect 496353 604208 500960 604210
rect 496353 604152 496358 604208
rect 496414 604152 500960 604208
rect 496353 604150 500960 604152
rect 496353 604147 496419 604150
rect 499520 604060 500960 604150
rect -960 599858 480 599948
rect 3509 599858 3575 599861
rect -960 599856 3575 599858
rect -960 599800 3514 599856
rect 3570 599800 3575 599856
rect -960 599798 3575 599800
rect -960 599708 480 599798
rect 3509 599795 3575 599798
rect 495433 599586 495499 599589
rect 499520 599586 500960 599676
rect 495433 599584 500960 599586
rect 495433 599528 495438 599584
rect 495494 599528 500960 599584
rect 495433 599526 500960 599528
rect 495433 599523 495499 599526
rect 499520 599436 500960 599526
rect 50153 599042 50219 599045
rect 50286 599042 50292 599044
rect 50153 599040 50292 599042
rect 50153 598984 50158 599040
rect 50214 598984 50292 599040
rect 50153 598982 50292 598984
rect 50153 598979 50219 598982
rect 50286 598980 50292 598982
rect 50356 598980 50362 599044
rect 70894 596396 70900 596460
rect 70964 596458 70970 596460
rect 205449 596458 205515 596461
rect 70964 596456 205515 596458
rect 70964 596400 205454 596456
rect 205510 596400 205515 596456
rect 70964 596398 205515 596400
rect 70964 596396 70970 596398
rect 205449 596395 205515 596398
rect 205909 596324 205975 596325
rect 205909 596320 205956 596324
rect 206020 596322 206026 596324
rect 205909 596264 205914 596320
rect 205909 596260 205956 596264
rect 206020 596262 206066 596322
rect 206020 596260 206026 596262
rect 205909 596259 205975 596260
rect -960 595506 480 595596
rect 2773 595506 2839 595509
rect -960 595504 2839 595506
rect -960 595448 2778 595504
rect 2834 595448 2839 595504
rect -960 595446 2839 595448
rect -960 595356 480 595446
rect 2773 595443 2839 595446
rect 496261 595234 496327 595237
rect 499520 595234 500960 595324
rect 496261 595232 500960 595234
rect 496261 595176 496266 595232
rect 496322 595176 500960 595232
rect 496261 595174 500960 595176
rect 496261 595171 496327 595174
rect 499520 595084 500960 595174
rect -960 590732 480 590972
rect 499520 590732 500960 590972
rect -960 586530 480 586620
rect 2773 586530 2839 586533
rect -960 586470 1042 586530
rect -960 586380 480 586470
rect 982 586394 1042 586470
rect 2638 586528 2839 586530
rect 2638 586472 2778 586528
rect 2834 586472 2839 586528
rect 2638 586470 2839 586472
rect 2638 586394 2698 586470
rect 2773 586467 2839 586470
rect 982 586334 2698 586394
rect 499520 586108 500960 586348
rect 201493 583812 201559 583813
rect 201493 583808 201540 583812
rect 201604 583810 201610 583812
rect 201493 583752 201498 583808
rect 201493 583748 201540 583752
rect 201604 583750 201650 583810
rect 201604 583748 201610 583750
rect 201493 583747 201559 583748
rect -960 581756 480 581996
rect 499520 581756 500960 581996
rect -960 577554 480 577644
rect 2773 577554 2839 577557
rect -960 577552 2839 577554
rect -960 577496 2778 577552
rect 2834 577496 2839 577552
rect -960 577494 2839 577496
rect -960 577404 480 577494
rect 2773 577491 2839 577494
rect 499520 577132 500960 577372
rect -960 573052 480 573292
rect 495433 572930 495499 572933
rect 499520 572930 500960 573020
rect 495433 572928 500960 572930
rect 495433 572872 495438 572928
rect 495494 572872 500960 572928
rect 495433 572870 500960 572872
rect 495433 572867 495499 572870
rect 499520 572780 500960 572870
rect -960 568428 480 568668
rect 499520 568156 500960 568396
rect 75913 566130 75979 566133
rect 111006 566130 111012 566132
rect 75913 566128 111012 566130
rect 75913 566072 75918 566128
rect 75974 566072 111012 566128
rect 75913 566070 111012 566072
rect 75913 566067 75979 566070
rect 111006 566068 111012 566070
rect 111076 566068 111082 566132
rect 76281 565858 76347 565861
rect 76414 565858 76420 565860
rect 76281 565856 76420 565858
rect 76281 565800 76286 565856
rect 76342 565800 76420 565856
rect 76281 565798 76420 565800
rect 76281 565795 76347 565798
rect 76414 565796 76420 565798
rect 76484 565796 76490 565860
rect -960 564076 480 564316
rect 499520 563804 500960 564044
rect -960 559602 480 559692
rect 2865 559602 2931 559605
rect -960 559600 2931 559602
rect -960 559544 2870 559600
rect 2926 559544 2931 559600
rect -960 559542 2931 559544
rect -960 559452 480 559542
rect 2865 559539 2931 559542
rect 499520 559180 500960 559420
rect -960 555250 480 555340
rect 2773 555250 2839 555253
rect -960 555248 2839 555250
rect -960 555192 2778 555248
rect 2834 555192 2839 555248
rect -960 555190 2839 555192
rect -960 555100 480 555190
rect 2773 555187 2839 555190
rect 495433 554978 495499 554981
rect 499520 554978 500960 555068
rect 495433 554976 500960 554978
rect 495433 554920 495438 554976
rect 495494 554920 500960 554976
rect 495433 554918 500960 554920
rect 495433 554915 495499 554918
rect 499520 554828 500960 554918
rect 268285 553484 268351 553485
rect 268285 553480 268332 553484
rect 268396 553482 268402 553484
rect 268561 553482 268627 553485
rect 276606 553482 276612 553484
rect 268285 553424 268290 553480
rect 268285 553420 268332 553424
rect 268396 553422 268442 553482
rect 268561 553480 276612 553482
rect 268561 553424 268566 553480
rect 268622 553424 276612 553480
rect 268561 553422 276612 553424
rect 268396 553420 268402 553422
rect 268285 553419 268351 553420
rect 268561 553419 268627 553422
rect 276606 553420 276612 553422
rect 276676 553420 276682 553484
rect -960 550476 480 550716
rect 495433 550354 495499 550357
rect 499520 550354 500960 550444
rect 495433 550352 500960 550354
rect 495433 550296 495438 550352
rect 495494 550296 500960 550352
rect 495433 550294 500960 550296
rect 495433 550291 495499 550294
rect 499520 550204 500960 550294
rect -960 546274 480 546364
rect 3141 546274 3207 546277
rect -960 546272 3207 546274
rect -960 546216 3146 546272
rect 3202 546216 3207 546272
rect -960 546214 3207 546216
rect -960 546124 480 546214
rect 3141 546211 3207 546214
rect 495433 546002 495499 546005
rect 499520 546002 500960 546092
rect 495433 546000 500960 546002
rect 495433 545944 495438 546000
rect 495494 545944 500960 546000
rect 495433 545942 500960 545944
rect 495433 545939 495499 545942
rect 499520 545852 500960 545942
rect 157425 543826 157491 543829
rect 157558 543826 157564 543828
rect 157425 543824 157564 543826
rect 157425 543768 157430 543824
rect 157486 543768 157564 543824
rect 157425 543766 157564 543768
rect 157425 543763 157491 543766
rect 157558 543764 157564 543766
rect 157628 543764 157634 543828
rect -960 541650 480 541740
rect 2865 541650 2931 541653
rect -960 541648 2931 541650
rect -960 541592 2870 541648
rect 2926 541592 2931 541648
rect -960 541590 2931 541592
rect -960 541500 480 541590
rect 2865 541587 2931 541590
rect 123293 541652 123359 541653
rect 123293 541648 123340 541652
rect 123404 541650 123410 541652
rect 123293 541592 123298 541648
rect 123293 541588 123340 541592
rect 123404 541590 123450 541650
rect 123404 541588 123410 541590
rect 123293 541587 123359 541588
rect 119981 541514 120047 541517
rect 128854 541514 128860 541516
rect 119981 541512 128860 541514
rect 119981 541456 119986 541512
rect 120042 541456 128860 541512
rect 119981 541454 128860 541456
rect 119981 541451 120047 541454
rect 128854 541452 128860 541454
rect 128924 541452 128930 541516
rect 495433 541378 495499 541381
rect 499520 541378 500960 541468
rect 495433 541376 500960 541378
rect 495433 541320 495438 541376
rect 495494 541320 500960 541376
rect 495433 541318 500960 541320
rect 495433 541315 495499 541318
rect 499520 541228 500960 541318
rect 159081 539610 159147 539613
rect 159214 539610 159220 539612
rect 159081 539608 159220 539610
rect 159081 539552 159086 539608
rect 159142 539552 159220 539608
rect 159081 539550 159220 539552
rect 159081 539547 159147 539550
rect 159214 539548 159220 539550
rect 159284 539548 159290 539612
rect -960 537298 480 537388
rect 3141 537298 3207 537301
rect -960 537296 3207 537298
rect -960 537240 3146 537296
rect 3202 537240 3207 537296
rect -960 537238 3207 537240
rect -960 537148 480 537238
rect 3141 537235 3207 537238
rect 495433 537026 495499 537029
rect 499520 537026 500960 537116
rect 495433 537024 500960 537026
rect 495433 536968 495438 537024
rect 495494 536968 500960 537024
rect 495433 536966 500960 536968
rect 495433 536963 495499 536966
rect 499520 536876 500960 536966
rect -960 532524 480 532764
rect 496077 532674 496143 532677
rect 499520 532674 500960 532764
rect 496077 532672 500960 532674
rect 496077 532616 496082 532672
rect 496138 532616 500960 532672
rect 496077 532614 500960 532616
rect 496077 532611 496143 532614
rect 499520 532524 500960 532614
rect -960 528322 480 528412
rect 3693 528322 3759 528325
rect -960 528320 3759 528322
rect -960 528264 3698 528320
rect 3754 528264 3759 528320
rect -960 528262 3759 528264
rect -960 528172 480 528262
rect 3693 528259 3759 528262
rect 495433 528050 495499 528053
rect 499520 528050 500960 528140
rect 495433 528048 500960 528050
rect 495433 527992 495438 528048
rect 495494 527992 500960 528048
rect 495433 527990 500960 527992
rect 495433 527987 495499 527990
rect 499520 527900 500960 527990
rect 117078 525268 117084 525332
rect 117148 525330 117154 525332
rect 262765 525330 262831 525333
rect 117148 525328 262831 525330
rect 117148 525272 262770 525328
rect 262826 525272 262831 525328
rect 117148 525270 262831 525272
rect 117148 525268 117154 525270
rect 262765 525267 262831 525270
rect 139894 525132 139900 525196
rect 139964 525194 139970 525196
rect 262673 525194 262739 525197
rect 139964 525192 262739 525194
rect 139964 525136 262678 525192
rect 262734 525136 262739 525192
rect 139964 525134 262739 525136
rect 139964 525132 139970 525134
rect 262673 525131 262739 525134
rect -960 523548 480 523788
rect 499520 523548 500960 523788
rect -960 519346 480 519436
rect 3877 519346 3943 519349
rect -960 519344 3943 519346
rect -960 519288 3882 519344
rect 3938 519288 3943 519344
rect -960 519286 3943 519288
rect -960 519196 480 519286
rect 3877 519283 3943 519286
rect 499520 518924 500960 519164
rect 96470 518740 96476 518804
rect 96540 518802 96546 518804
rect 291101 518802 291167 518805
rect 96540 518800 291167 518802
rect 96540 518744 291106 518800
rect 291162 518744 291167 518800
rect 96540 518742 291167 518744
rect 96540 518740 96546 518742
rect 291101 518739 291167 518742
rect 112294 518604 112300 518668
rect 112364 518666 112370 518668
rect 289813 518666 289879 518669
rect 112364 518664 289879 518666
rect 112364 518608 289818 518664
rect 289874 518608 289879 518664
rect 112364 518606 289879 518608
rect 112364 518604 112370 518606
rect 289813 518603 289879 518606
rect -960 514994 480 515084
rect 3325 514994 3391 514997
rect -960 514992 3391 514994
rect -960 514936 3330 514992
rect 3386 514936 3391 514992
rect -960 514934 3391 514936
rect -960 514844 480 514934
rect 3325 514931 3391 514934
rect 499520 514572 500960 514812
rect -960 510220 480 510460
rect 495433 510098 495499 510101
rect 499520 510098 500960 510188
rect 495433 510096 500960 510098
rect 495433 510040 495438 510096
rect 495494 510040 500960 510096
rect 495433 510038 500960 510040
rect 495433 510035 495499 510038
rect 499520 509948 500960 510038
rect -960 506018 480 506108
rect 3141 506018 3207 506021
rect -960 506016 3207 506018
rect -960 505960 3146 506016
rect 3202 505960 3207 506016
rect -960 505958 3207 505960
rect -960 505868 480 505958
rect 3141 505955 3207 505958
rect 499520 505596 500960 505836
rect -960 501244 480 501484
rect 499520 500972 500960 501212
rect 190361 499628 190427 499629
rect 190310 499626 190316 499628
rect 190270 499566 190316 499626
rect 190380 499624 190427 499628
rect 190422 499568 190427 499624
rect 190310 499564 190316 499566
rect 190380 499564 190427 499568
rect 190361 499563 190427 499564
rect 208577 498130 208643 498133
rect 220854 498130 220860 498132
rect 208577 498128 220860 498130
rect 208577 498072 208582 498128
rect 208638 498072 220860 498128
rect 208577 498070 220860 498072
rect 208577 498067 208643 498070
rect 220854 498068 220860 498070
rect 220924 498068 220930 498132
rect -960 497042 480 497132
rect 2773 497042 2839 497045
rect -960 497040 2839 497042
rect -960 496984 2778 497040
rect 2834 496984 2839 497040
rect -960 496982 2839 496984
rect -960 496892 480 496982
rect 2773 496979 2839 496982
rect 499520 496620 500960 496860
rect 32305 493098 32371 493101
rect 57094 493098 57100 493100
rect 32305 493096 57100 493098
rect 32305 493040 32310 493096
rect 32366 493040 57100 493096
rect 32305 493038 57100 493040
rect 32305 493035 32371 493038
rect 57094 493036 57100 493038
rect 57164 493036 57170 493100
rect 32397 492692 32463 492693
rect 32397 492688 32444 492692
rect 32508 492690 32514 492692
rect 32397 492632 32402 492688
rect 32397 492628 32444 492632
rect 32508 492630 32554 492690
rect 32508 492628 32514 492630
rect 32397 492627 32463 492628
rect -960 492268 480 492508
rect 499520 491996 500960 492236
rect -960 487916 480 488156
rect 499520 487644 500960 487884
rect -960 483292 480 483532
rect 499520 483020 500960 483260
rect -960 479090 480 479180
rect 2773 479090 2839 479093
rect -960 479088 2839 479090
rect -960 479032 2778 479088
rect 2834 479032 2839 479088
rect -960 479030 2839 479032
rect -960 478940 480 479030
rect 2773 479027 2839 479030
rect 496353 478818 496419 478821
rect 499520 478818 500960 478908
rect 496353 478816 500960 478818
rect 496353 478760 496358 478816
rect 496414 478760 500960 478816
rect 496353 478758 500960 478760
rect 496353 478755 496419 478758
rect 499520 478668 500960 478758
rect -960 474316 480 474556
rect 496445 474466 496511 474469
rect 499520 474466 500960 474556
rect 496445 474464 500960 474466
rect 496445 474408 496450 474464
rect 496506 474408 500960 474464
rect 496445 474406 500960 474408
rect 496445 474403 496511 474406
rect 499520 474316 500960 474406
rect 93761 473514 93827 473517
rect 145414 473514 145420 473516
rect 93761 473512 145420 473514
rect 93761 473456 93766 473512
rect 93822 473456 145420 473512
rect 93761 473454 145420 473456
rect 93761 473451 93827 473454
rect 145414 473452 145420 473454
rect 145484 473452 145490 473516
rect 198273 470658 198339 470661
rect 200614 470658 200620 470660
rect 198273 470656 200620 470658
rect 198273 470600 198278 470656
rect 198334 470600 200620 470656
rect 198273 470598 200620 470600
rect 198273 470595 198339 470598
rect 200614 470596 200620 470598
rect 200684 470596 200690 470660
rect -960 469964 480 470204
rect 495433 469842 495499 469845
rect 499520 469842 500960 469932
rect 495433 469840 500960 469842
rect 495433 469784 495438 469840
rect 495494 469784 500960 469840
rect 495433 469782 500960 469784
rect 495433 469779 495499 469782
rect 499520 469692 500960 469782
rect -960 465340 480 465580
rect 499520 465340 500960 465580
rect -960 461138 480 461228
rect 3325 461138 3391 461141
rect -960 461136 3391 461138
rect -960 461080 3330 461136
rect 3386 461080 3391 461136
rect -960 461078 3391 461080
rect -960 460988 480 461078
rect 3325 461075 3391 461078
rect 499520 460716 500960 460956
rect -960 456636 480 456876
rect 495433 456514 495499 456517
rect 499520 456514 500960 456604
rect 495433 456512 500960 456514
rect 495433 456456 495438 456512
rect 495494 456456 500960 456512
rect 495433 456454 500960 456456
rect 495433 456451 495499 456454
rect 499520 456364 500960 456454
rect -960 452012 480 452252
rect 496537 451890 496603 451893
rect 499520 451890 500960 451980
rect 496537 451888 500960 451890
rect 496537 451832 496542 451888
rect 496598 451832 500960 451888
rect 496537 451830 500960 451832
rect 496537 451827 496603 451830
rect 499520 451740 500960 451830
rect -960 447660 480 447900
rect 499520 447388 500960 447628
rect 112345 446994 112411 446997
rect 146886 446994 146892 446996
rect 112345 446992 146892 446994
rect 112345 446936 112350 446992
rect 112406 446936 146892 446992
rect 112345 446934 146892 446936
rect 112345 446931 112411 446934
rect 146886 446932 146892 446934
rect 146956 446932 146962 446996
rect -960 443186 480 443276
rect 3141 443186 3207 443189
rect -960 443184 3207 443186
rect -960 443128 3146 443184
rect 3202 443128 3207 443184
rect -960 443126 3207 443128
rect -960 443036 480 443126
rect 3141 443123 3207 443126
rect 152365 443050 152431 443053
rect 155166 443050 155172 443052
rect 152365 443048 155172 443050
rect 152365 442992 152370 443048
rect 152426 442992 155172 443048
rect 152365 442990 155172 442992
rect 152365 442987 152431 442990
rect 155166 442988 155172 442990
rect 155236 442988 155242 443052
rect 495433 442914 495499 442917
rect 499520 442914 500960 443004
rect 495433 442912 500960 442914
rect 495433 442856 495438 442912
rect 495494 442856 500960 442912
rect 495433 442854 500960 442856
rect 495433 442851 495499 442854
rect 499520 442764 500960 442854
rect -960 438684 480 438924
rect 499520 438412 500960 438652
rect 263685 436116 263751 436117
rect 263685 436112 263732 436116
rect 263796 436114 263802 436116
rect 263685 436056 263690 436112
rect 263685 436052 263732 436056
rect 263796 436054 263842 436114
rect 263796 436052 263802 436054
rect 263685 436051 263751 436052
rect 34278 434964 34284 435028
rect 34348 435026 34354 435028
rect 47669 435026 47735 435029
rect 34348 435024 47735 435026
rect 34348 434968 47674 435024
rect 47730 434968 47735 435024
rect 34348 434966 47735 434968
rect 34348 434964 34354 434966
rect 47669 434963 47735 434966
rect 48037 434756 48103 434757
rect 48037 434752 48084 434756
rect 48148 434754 48154 434756
rect 48037 434696 48042 434752
rect 48037 434692 48084 434696
rect 48148 434694 48194 434754
rect 48148 434692 48154 434694
rect 48037 434691 48103 434692
rect -960 434210 480 434300
rect 3325 434210 3391 434213
rect -960 434208 3391 434210
rect -960 434152 3330 434208
rect 3386 434152 3391 434208
rect -960 434150 3391 434152
rect -960 434060 480 434150
rect 3325 434147 3391 434150
rect 499520 433788 500960 434028
rect 86166 433332 86172 433396
rect 86236 433394 86242 433396
rect 91461 433394 91527 433397
rect 86236 433392 91527 433394
rect 86236 433336 91466 433392
rect 91522 433336 91527 433392
rect 86236 433334 91527 433336
rect 86236 433332 86242 433334
rect 91461 433331 91527 433334
rect 36486 432108 36492 432172
rect 36556 432170 36562 432172
rect 281625 432170 281691 432173
rect 36556 432168 281691 432170
rect 36556 432112 281630 432168
rect 281686 432112 281691 432168
rect 36556 432110 281691 432112
rect 36556 432108 36562 432110
rect 281625 432107 281691 432110
rect 282729 432036 282795 432037
rect 282678 432034 282684 432036
rect 282638 431974 282684 432034
rect 282748 432032 282795 432036
rect 282790 431976 282795 432032
rect 282678 431972 282684 431974
rect 282748 431972 282795 431976
rect 282729 431971 282795 431972
rect -960 429858 480 429948
rect 3233 429858 3299 429861
rect -960 429856 3299 429858
rect -960 429800 3238 429856
rect 3294 429800 3299 429856
rect -960 429798 3299 429800
rect -960 429708 480 429798
rect 3233 429795 3299 429798
rect 499520 429436 500960 429676
rect -960 425234 480 425324
rect 3325 425234 3391 425237
rect -960 425232 3391 425234
rect -960 425176 3330 425232
rect 3386 425176 3391 425232
rect -960 425174 3391 425176
rect -960 425084 480 425174
rect 3325 425171 3391 425174
rect 499520 424812 500960 425052
rect -960 420882 480 420972
rect 3693 420882 3759 420885
rect -960 420880 3759 420882
rect -960 420824 3698 420880
rect 3754 420824 3759 420880
rect -960 420822 3759 420824
rect -960 420732 480 420822
rect 3693 420819 3759 420822
rect 495985 420610 496051 420613
rect 499520 420610 500960 420700
rect 495985 420608 500960 420610
rect 495985 420552 495990 420608
rect 496046 420552 500960 420608
rect 495985 420550 500960 420552
rect 495985 420547 496051 420550
rect 499520 420460 500960 420550
rect -960 416258 480 416348
rect 3785 416258 3851 416261
rect -960 416256 3851 416258
rect -960 416200 3790 416256
rect 3846 416200 3851 416256
rect -960 416198 3851 416200
rect -960 416108 480 416198
rect 3785 416195 3851 416198
rect 499520 416108 500960 416348
rect 119613 414084 119679 414085
rect 119613 414080 119660 414084
rect 119724 414082 119730 414084
rect 119613 414024 119618 414080
rect 119613 414020 119660 414024
rect 119724 414022 119770 414082
rect 119724 414020 119730 414022
rect 119613 414019 119679 414020
rect -960 411756 480 411996
rect 499520 411484 500960 411724
rect 48814 410484 48820 410548
rect 48884 410546 48890 410548
rect 112805 410546 112871 410549
rect 48884 410544 112871 410546
rect 48884 410488 112810 410544
rect 112866 410488 112871 410544
rect 48884 410486 112871 410488
rect 48884 410484 48890 410486
rect 112805 410483 112871 410486
rect 55305 410002 55371 410005
rect 55438 410002 55444 410004
rect 55305 410000 55444 410002
rect 55305 409944 55310 410000
rect 55366 409944 55444 410000
rect 55305 409942 55444 409944
rect 55305 409939 55371 409942
rect 55438 409940 55444 409942
rect 55508 409940 55514 410004
rect -960 407282 480 407372
rect 3325 407282 3391 407285
rect -960 407280 3391 407282
rect -960 407224 3330 407280
rect 3386 407224 3391 407280
rect -960 407222 3391 407224
rect -960 407132 480 407222
rect 3325 407219 3391 407222
rect 495433 407282 495499 407285
rect 499520 407282 500960 407372
rect 495433 407280 500960 407282
rect 495433 407224 495438 407280
rect 495494 407224 500960 407280
rect 495433 407222 500960 407224
rect 495433 407219 495499 407222
rect 499520 407132 500960 407222
rect -960 402930 480 403020
rect 2957 402930 3023 402933
rect -960 402928 3023 402930
rect -960 402872 2962 402928
rect 3018 402872 3023 402928
rect -960 402870 3023 402872
rect -960 402780 480 402870
rect 2957 402867 3023 402870
rect 495433 402658 495499 402661
rect 499520 402658 500960 402748
rect 495433 402656 500960 402658
rect 495433 402600 495438 402656
rect 495494 402600 500960 402656
rect 495433 402598 500960 402600
rect 495433 402595 495499 402598
rect 499520 402508 500960 402598
rect 67357 400620 67423 400621
rect 67357 400618 67404 400620
rect 67312 400616 67404 400618
rect 67468 400618 67474 400620
rect 67541 400618 67607 400621
rect 67468 400616 67607 400618
rect 67312 400560 67362 400616
rect 67468 400560 67546 400616
rect 67602 400560 67607 400616
rect 67312 400558 67404 400560
rect 67357 400556 67404 400558
rect 67468 400558 67607 400560
rect 67468 400556 67474 400558
rect 67357 400555 67423 400556
rect 67541 400555 67607 400558
rect 67633 400346 67699 400349
rect 69606 400346 69612 400348
rect 67633 400344 69612 400346
rect 67633 400288 67638 400344
rect 67694 400288 69612 400344
rect 67633 400286 69612 400288
rect 67633 400283 67699 400286
rect 69606 400284 69612 400286
rect 69676 400284 69682 400348
rect -960 398428 480 398668
rect 495433 398306 495499 398309
rect 499520 398306 500960 398396
rect 495433 398304 500960 398306
rect 495433 398248 495438 398304
rect 495494 398248 500960 398304
rect 495433 398246 500960 398248
rect 495433 398243 495499 398246
rect 499520 398156 500960 398246
rect -960 393804 480 394044
rect 499520 393532 500960 393772
rect -960 389602 480 389692
rect 3601 389602 3667 389605
rect -960 389600 3667 389602
rect -960 389544 3606 389600
rect 3662 389544 3667 389600
rect -960 389542 3667 389544
rect -960 389452 480 389542
rect 3601 389539 3667 389542
rect 499520 389180 500960 389420
rect -960 384978 480 385068
rect 3785 384978 3851 384981
rect -960 384976 3851 384978
rect -960 384920 3790 384976
rect 3846 384920 3851 384976
rect -960 384918 3851 384920
rect -960 384828 480 384918
rect 3785 384915 3851 384918
rect 495433 384706 495499 384709
rect 499520 384706 500960 384796
rect 495433 384704 500960 384706
rect 495433 384648 495438 384704
rect 495494 384648 500960 384704
rect 495433 384646 500960 384648
rect 495433 384643 495499 384646
rect 499520 384556 500960 384646
rect 132585 384298 132651 384301
rect 132718 384298 132724 384300
rect 132585 384296 132724 384298
rect 132585 384240 132590 384296
rect 132646 384240 132724 384296
rect 132585 384238 132724 384240
rect 132585 384235 132651 384238
rect 132718 384236 132724 384238
rect 132788 384236 132794 384300
rect 103513 384162 103579 384165
rect 103646 384162 103652 384164
rect 103513 384160 103652 384162
rect 103513 384104 103518 384160
rect 103574 384104 103652 384160
rect 103513 384102 103652 384104
rect 103513 384099 103579 384102
rect 103646 384100 103652 384102
rect 103716 384100 103722 384164
rect 88793 384026 88859 384029
rect 88926 384026 88932 384028
rect 88793 384024 88932 384026
rect 88793 383968 88798 384024
rect 88854 383968 88932 384024
rect 88793 383966 88932 383968
rect 88793 383963 88859 383966
rect 88926 383964 88932 383966
rect 88996 383964 89002 384028
rect 37774 383828 37780 383892
rect 37844 383890 37850 383892
rect 177205 383890 177271 383893
rect 37844 383888 177271 383890
rect 37844 383832 177210 383888
rect 177266 383832 177271 383888
rect 37844 383830 177271 383832
rect 37844 383828 37850 383830
rect 177205 383827 177271 383830
rect 38878 380972 38884 381036
rect 38948 381034 38954 381036
rect 39389 381034 39455 381037
rect 38948 381032 39455 381034
rect 38948 380976 39394 381032
rect 39450 380976 39455 381032
rect 38948 380974 39455 380976
rect 38948 380972 38954 380974
rect 39389 380971 39455 380974
rect -960 380476 480 380716
rect 72918 380428 72924 380492
rect 72988 380490 72994 380492
rect 274449 380490 274515 380493
rect 72988 380488 274515 380490
rect 72988 380432 274454 380488
rect 274510 380432 274515 380488
rect 72988 380430 274515 380432
rect 72988 380428 72994 380430
rect 274449 380427 274515 380430
rect 499520 380204 500960 380444
rect -960 375852 480 376092
rect 499520 375580 500960 375820
rect 233693 371788 233759 371789
rect 233693 371786 233740 371788
rect 233648 371784 233740 371786
rect -960 371500 480 371740
rect 233648 371728 233698 371784
rect 233648 371726 233740 371728
rect 233693 371724 233740 371726
rect 233804 371724 233810 371788
rect 233693 371723 233759 371724
rect 499520 371228 500960 371468
rect 214741 369882 214807 369885
rect 217174 369882 217180 369884
rect 214741 369880 217180 369882
rect 214741 369824 214746 369880
rect 214802 369824 217180 369880
rect 214741 369822 217180 369824
rect 214741 369819 214807 369822
rect 217174 369820 217180 369822
rect 217244 369820 217250 369884
rect -960 367026 480 367116
rect 2773 367026 2839 367029
rect -960 367024 2839 367026
rect -960 366968 2778 367024
rect 2834 366968 2839 367024
rect -960 366966 2839 366968
rect -960 366876 480 366966
rect 2773 366963 2839 366966
rect 495433 366754 495499 366757
rect 499520 366754 500960 366844
rect 495433 366752 500960 366754
rect 495433 366696 495438 366752
rect 495494 366696 500960 366752
rect 495433 366694 500960 366696
rect 495433 366691 495499 366694
rect 499520 366604 500960 366694
rect 143073 365394 143139 365397
rect 143206 365394 143212 365396
rect 143073 365392 143212 365394
rect 143073 365336 143078 365392
rect 143134 365336 143212 365392
rect 143073 365334 143212 365336
rect 143073 365331 143139 365334
rect 143206 365332 143212 365334
rect 143276 365332 143282 365396
rect -960 362524 480 362764
rect 180057 362538 180123 362541
rect 196566 362538 196572 362540
rect 180057 362536 196572 362538
rect 180057 362480 180062 362536
rect 180118 362480 196572 362536
rect 180057 362478 196572 362480
rect 180057 362475 180123 362478
rect 196566 362476 196572 362478
rect 196636 362476 196642 362540
rect 495433 362402 495499 362405
rect 499520 362402 500960 362492
rect 495433 362400 500960 362402
rect 495433 362344 495438 362400
rect 495494 362344 500960 362400
rect 495433 362342 500960 362344
rect 495433 362339 495499 362342
rect 499520 362252 500960 362342
rect -960 357900 480 358140
rect 496353 358050 496419 358053
rect 499520 358050 500960 358140
rect 496353 358048 500960 358050
rect 496353 357992 496358 358048
rect 496414 357992 500960 358048
rect 496353 357990 500960 357992
rect 496353 357987 496419 357990
rect 499520 357900 500960 357990
rect 90633 356554 90699 356557
rect 99414 356554 99420 356556
rect 90633 356552 99420 356554
rect 90633 356496 90638 356552
rect 90694 356496 99420 356552
rect 90633 356494 99420 356496
rect 90633 356491 90699 356494
rect 99414 356492 99420 356494
rect 99484 356492 99490 356556
rect -960 353548 480 353788
rect 117814 353364 117820 353428
rect 117884 353426 117890 353428
rect 194593 353426 194659 353429
rect 117884 353424 194659 353426
rect 117884 353368 194598 353424
rect 194654 353368 194659 353424
rect 117884 353366 194659 353368
rect 117884 353364 117890 353366
rect 194593 353363 194659 353366
rect 499520 353276 500960 353516
rect -960 348924 480 349164
rect 499520 348924 500960 349164
rect -960 344572 480 344812
rect 499520 344300 500960 344540
rect -960 340220 480 340460
rect 499520 339948 500960 340188
rect 218697 337650 218763 337653
rect 223614 337650 223620 337652
rect 218697 337648 223620 337650
rect 218697 337592 218702 337648
rect 218758 337592 223620 337648
rect 218697 337590 223620 337592
rect 218697 337587 218763 337590
rect 223614 337588 223620 337590
rect 223684 337588 223690 337652
rect 231025 337380 231091 337381
rect 230974 337378 230980 337380
rect 230934 337318 230980 337378
rect 231044 337376 231091 337380
rect 231086 337320 231091 337376
rect 230974 337316 230980 337318
rect 231044 337316 231091 337320
rect 231025 337315 231091 337316
rect -960 335596 480 335836
rect 499520 335324 500960 335564
rect 38837 333300 38903 333301
rect 38837 333298 38884 333300
rect 38792 333296 38884 333298
rect 38792 333240 38842 333296
rect 38792 333238 38884 333240
rect 38837 333236 38884 333238
rect 38948 333236 38954 333300
rect 38837 333235 38903 333236
rect -960 331394 480 331484
rect 3601 331394 3667 331397
rect -960 331392 3667 331394
rect -960 331336 3606 331392
rect 3662 331336 3667 331392
rect -960 331334 3667 331336
rect -960 331244 480 331334
rect 3601 331331 3667 331334
rect 499520 330972 500960 331212
rect -960 326620 480 326860
rect 499520 326348 500960 326588
rect 263358 324940 263364 325004
rect 263428 325002 263434 325004
rect 282269 325002 282335 325005
rect 263428 325000 282335 325002
rect 263428 324944 282274 325000
rect 282330 324944 282335 325000
rect 263428 324942 282335 324944
rect 263428 324940 263434 324942
rect 282269 324939 282335 324942
rect -960 322418 480 322508
rect 3601 322418 3667 322421
rect -960 322416 3667 322418
rect -960 322360 3606 322416
rect 3662 322360 3667 322416
rect -960 322358 3667 322360
rect -960 322268 480 322358
rect 3601 322355 3667 322358
rect 495433 322146 495499 322149
rect 499520 322146 500960 322236
rect 495433 322144 500960 322146
rect 495433 322088 495438 322144
rect 495494 322088 500960 322144
rect 495433 322086 500960 322088
rect 495433 322083 495499 322086
rect 499520 321996 500960 322086
rect -960 317794 480 317884
rect 3049 317794 3115 317797
rect -960 317792 3115 317794
rect -960 317736 3054 317792
rect 3110 317736 3115 317792
rect -960 317734 3115 317736
rect -960 317644 480 317734
rect 3049 317731 3115 317734
rect 499520 317372 500960 317612
rect -960 313292 480 313532
rect 495433 313170 495499 313173
rect 499520 313170 500960 313260
rect 495433 313168 500960 313170
rect 495433 313112 495438 313168
rect 495494 313112 500960 313168
rect 495433 313110 500960 313112
rect 495433 313107 495499 313110
rect 499520 313020 500960 313110
rect -960 308818 480 308908
rect 4153 308818 4219 308821
rect -960 308816 4219 308818
rect -960 308760 4158 308816
rect 4214 308760 4219 308816
rect -960 308758 4219 308760
rect -960 308668 480 308758
rect 4153 308755 4219 308758
rect 495433 308546 495499 308549
rect 499520 308546 500960 308636
rect 495433 308544 500960 308546
rect 495433 308488 495438 308544
rect 495494 308488 500960 308544
rect 495433 308486 500960 308488
rect 495433 308483 495499 308486
rect 499520 308396 500960 308486
rect 140773 307050 140839 307053
rect 149646 307050 149652 307052
rect 140773 307048 149652 307050
rect 140773 306992 140778 307048
rect 140834 306992 149652 307048
rect 140773 306990 149652 306992
rect 140773 306987 140839 306990
rect 149646 306988 149652 306990
rect 149716 306988 149722 307052
rect -960 304316 480 304556
rect 499520 304044 500960 304284
rect 261109 300932 261175 300933
rect 261109 300928 261156 300932
rect 261220 300930 261226 300932
rect 261109 300872 261114 300928
rect 261109 300868 261156 300872
rect 261220 300870 261266 300930
rect 261220 300868 261226 300870
rect 261109 300867 261175 300868
rect -960 299692 480 299932
rect 495433 299842 495499 299845
rect 499520 299842 500960 299932
rect 495433 299840 500960 299842
rect 495433 299784 495438 299840
rect 495494 299784 500960 299840
rect 495433 299782 500960 299784
rect 495433 299779 495499 299782
rect 499520 299692 500960 299782
rect 112161 295626 112227 295629
rect 113766 295626 113772 295628
rect 112161 295624 113772 295626
rect -960 295340 480 295580
rect 112161 295568 112166 295624
rect 112222 295568 113772 295624
rect 112161 295566 113772 295568
rect 112161 295563 112227 295566
rect 113766 295564 113772 295566
rect 113836 295626 113842 295628
rect 114461 295626 114527 295629
rect 113836 295624 114527 295626
rect 113836 295568 114466 295624
rect 114522 295568 114527 295624
rect 113836 295566 114527 295568
rect 113836 295564 113842 295566
rect 114461 295563 114527 295566
rect 495433 295218 495499 295221
rect 499520 295218 500960 295308
rect 495433 295216 500960 295218
rect 495433 295160 495438 295216
rect 495494 295160 500960 295216
rect 495433 295158 500960 295160
rect 495433 295155 495499 295158
rect 499520 295068 500960 295158
rect -960 290866 480 290956
rect 3601 290866 3667 290869
rect -960 290864 3667 290866
rect -960 290808 3606 290864
rect 3662 290808 3667 290864
rect -960 290806 3667 290808
rect -960 290716 480 290806
rect 3601 290803 3667 290806
rect 496629 290866 496695 290869
rect 499520 290866 500960 290956
rect 496629 290864 500960 290866
rect 496629 290808 496634 290864
rect 496690 290808 500960 290864
rect 496629 290806 500960 290808
rect 496629 290803 496695 290806
rect 499520 290716 500960 290806
rect 46054 288084 46060 288148
rect 46124 288146 46130 288148
rect 92933 288146 92999 288149
rect 46124 288144 92999 288146
rect 46124 288088 92938 288144
rect 92994 288088 92999 288144
rect 46124 288086 92999 288088
rect 46124 288084 46130 288086
rect 92933 288083 92999 288086
rect 93117 288146 93183 288149
rect 108246 288146 108252 288148
rect 93117 288144 108252 288146
rect 93117 288088 93122 288144
rect 93178 288088 108252 288144
rect 93117 288086 108252 288088
rect 93117 288083 93183 288086
rect 108246 288084 108252 288086
rect 108316 288084 108322 288148
rect 109534 286996 109540 287060
rect 109604 287058 109610 287060
rect 273621 287058 273687 287061
rect 109604 287056 273687 287058
rect 109604 287000 273626 287056
rect 273682 287000 273687 287056
rect 109604 286998 273687 287000
rect 109604 286996 109610 286998
rect 273621 286995 273687 286998
rect -960 286364 480 286604
rect 495433 286242 495499 286245
rect 499520 286242 500960 286332
rect 495433 286240 500960 286242
rect 495433 286184 495438 286240
rect 495494 286184 500960 286240
rect 495433 286182 500960 286184
rect 495433 286179 495499 286182
rect 499520 286092 500960 286182
rect 273989 285700 274055 285701
rect 273989 285698 274036 285700
rect 273944 285696 274036 285698
rect 273944 285640 273994 285696
rect 273944 285638 274036 285640
rect 273989 285636 274036 285638
rect 274100 285636 274106 285700
rect 273989 285635 274055 285636
rect -960 282012 480 282252
rect 495433 281890 495499 281893
rect 499520 281890 500960 281980
rect 495433 281888 500960 281890
rect 495433 281832 495438 281888
rect 495494 281832 500960 281888
rect 495433 281830 500960 281832
rect 495433 281827 495499 281830
rect 499520 281740 500960 281830
rect -960 277388 480 277628
rect 496261 277266 496327 277269
rect 499520 277266 500960 277356
rect 496261 277264 500960 277266
rect 496261 277208 496266 277264
rect 496322 277208 500960 277264
rect 496261 277206 500960 277208
rect 496261 277203 496327 277206
rect 499520 277116 500960 277206
rect 159265 273866 159331 273869
rect 248229 273868 248295 273869
rect 191046 273866 191052 273868
rect 159265 273864 191052 273866
rect 159265 273808 159270 273864
rect 159326 273808 191052 273864
rect 159265 273806 191052 273808
rect 159265 273803 159331 273806
rect 191046 273804 191052 273806
rect 191116 273804 191122 273868
rect 248229 273864 248276 273868
rect 248340 273866 248346 273868
rect 248229 273808 248234 273864
rect 248229 273804 248276 273808
rect 248340 273806 248386 273866
rect 248340 273804 248346 273806
rect 248229 273803 248295 273804
rect -960 273186 480 273276
rect 3601 273186 3667 273189
rect -960 273184 3667 273186
rect -960 273128 3606 273184
rect 3662 273128 3667 273184
rect -960 273126 3667 273128
rect -960 273036 480 273126
rect 3601 273123 3667 273126
rect 495985 272914 496051 272917
rect 499520 272914 500960 273004
rect 495985 272912 500960 272914
rect 495985 272856 495990 272912
rect 496046 272856 500960 272912
rect 495985 272854 500960 272856
rect 495985 272851 496051 272854
rect 499520 272764 500960 272854
rect -960 268562 480 268652
rect 3601 268562 3667 268565
rect -960 268560 3667 268562
rect -960 268504 3606 268560
rect 3662 268504 3667 268560
rect -960 268502 3667 268504
rect -960 268412 480 268502
rect 3601 268499 3667 268502
rect 495433 268290 495499 268293
rect 499520 268290 500960 268380
rect 495433 268288 500960 268290
rect 495433 268232 495438 268288
rect 495494 268232 500960 268288
rect 495433 268230 500960 268232
rect 495433 268227 495499 268230
rect 499520 268140 500960 268230
rect 216070 267820 216076 267884
rect 216140 267882 216146 267884
rect 229093 267882 229159 267885
rect 216140 267880 229159 267882
rect 216140 267824 229098 267880
rect 229154 267824 229159 267880
rect 216140 267822 229159 267824
rect 216140 267820 216146 267822
rect 229093 267819 229159 267822
rect 103421 266932 103487 266933
rect 103421 266930 103468 266932
rect 103376 266928 103468 266930
rect 103532 266930 103538 266932
rect 103376 266872 103426 266928
rect 103376 266870 103468 266872
rect 103421 266868 103468 266870
rect 103532 266870 103614 266930
rect 103532 266868 103538 266870
rect 103421 266867 103487 266868
rect -960 264210 480 264300
rect 3877 264210 3943 264213
rect -960 264208 3943 264210
rect -960 264152 3882 264208
rect 3938 264152 3943 264208
rect -960 264150 3943 264152
rect -960 264060 480 264150
rect 3877 264147 3943 264150
rect 499520 263788 500960 264028
rect 98729 263666 98795 263669
rect 98862 263666 98868 263668
rect 98729 263664 98868 263666
rect 98729 263608 98734 263664
rect 98790 263608 98868 263664
rect 98729 263606 98868 263608
rect 98729 263603 98795 263606
rect 98862 263604 98868 263606
rect 98932 263604 98938 263668
rect 207381 262444 207447 262445
rect 207381 262442 207428 262444
rect 207336 262440 207428 262442
rect 207336 262384 207386 262440
rect 207336 262382 207428 262384
rect 207381 262380 207428 262382
rect 207492 262380 207498 262444
rect 207381 262379 207447 262380
rect 125317 261218 125383 261221
rect 130326 261218 130332 261220
rect 125317 261216 130332 261218
rect 125317 261160 125322 261216
rect 125378 261160 130332 261216
rect 125317 261158 130332 261160
rect 125317 261155 125383 261158
rect 130326 261156 130332 261158
rect 130396 261218 130402 261220
rect 130469 261218 130535 261221
rect 130396 261216 130535 261218
rect 130396 261160 130474 261216
rect 130530 261160 130535 261216
rect 130396 261158 130535 261160
rect 130396 261156 130402 261158
rect 130469 261155 130535 261158
rect 125726 260884 125732 260948
rect 125796 260946 125802 260948
rect 125869 260946 125935 260949
rect 125796 260944 125935 260946
rect 125796 260888 125874 260944
rect 125930 260888 125935 260944
rect 125796 260886 125935 260888
rect 125796 260884 125802 260886
rect 125869 260883 125935 260886
rect 131573 260948 131639 260949
rect 131573 260944 131620 260948
rect 131684 260946 131690 260948
rect 131573 260888 131578 260944
rect 131573 260884 131620 260888
rect 131684 260886 131730 260946
rect 131684 260884 131690 260886
rect 131573 260883 131639 260884
rect -960 259436 480 259676
rect 495433 259314 495499 259317
rect 499520 259314 500960 259404
rect 495433 259312 500960 259314
rect 495433 259256 495438 259312
rect 495494 259256 500960 259312
rect 495433 259254 500960 259256
rect 495433 259251 495499 259254
rect 103278 259116 103284 259180
rect 103348 259178 103354 259180
rect 180885 259178 180951 259181
rect 103348 259176 180951 259178
rect 103348 259120 180890 259176
rect 180946 259120 180951 259176
rect 499520 259164 500960 259254
rect 103348 259118 180951 259120
rect 103348 259116 103354 259118
rect 180885 259115 180951 259118
rect 180793 258634 180859 258637
rect 180926 258634 180932 258636
rect 180793 258632 180932 258634
rect 180793 258576 180798 258632
rect 180854 258576 180932 258632
rect 180793 258574 180932 258576
rect 180793 258571 180859 258574
rect 180926 258572 180932 258574
rect 180996 258572 181002 258636
rect -960 255234 480 255324
rect 3877 255234 3943 255237
rect -960 255232 3943 255234
rect -960 255176 3882 255232
rect 3938 255176 3943 255232
rect -960 255174 3943 255176
rect -960 255084 480 255174
rect 3877 255171 3943 255174
rect 40534 254764 40540 254828
rect 40604 254826 40610 254828
rect 219801 254826 219867 254829
rect 40604 254824 219867 254826
rect 40604 254768 219806 254824
rect 219862 254768 219867 254824
rect 499520 254812 500960 255052
rect 40604 254766 219867 254768
rect 40604 254764 40610 254766
rect 219801 254763 219867 254766
rect 219249 254692 219315 254693
rect 219198 254628 219204 254692
rect 219268 254690 219315 254692
rect 219268 254688 219360 254690
rect 219310 254632 219360 254688
rect 219268 254630 219360 254632
rect 219268 254628 219315 254630
rect 219249 254627 219315 254628
rect -960 250460 480 250700
rect 495433 250338 495499 250341
rect 499520 250338 500960 250428
rect 495433 250336 500960 250338
rect 495433 250280 495438 250336
rect 495494 250280 500960 250336
rect 495433 250278 500960 250280
rect 495433 250275 495499 250278
rect 499520 250188 500960 250278
rect 303153 249930 303219 249933
rect 303286 249930 303292 249932
rect 303153 249928 303292 249930
rect 303153 249872 303158 249928
rect 303214 249872 303292 249928
rect 303153 249870 303292 249872
rect 303153 249867 303219 249870
rect 303286 249868 303292 249870
rect 303356 249868 303362 249932
rect 103421 248436 103487 248437
rect 103421 248434 103468 248436
rect 103376 248432 103468 248434
rect 103532 248434 103538 248436
rect 103376 248376 103426 248432
rect 103376 248374 103468 248376
rect 103421 248372 103468 248374
rect 103532 248374 103614 248434
rect 103532 248372 103538 248374
rect 103421 248371 103487 248372
rect -960 246258 480 246348
rect 3325 246258 3391 246261
rect -960 246256 3391 246258
rect -960 246200 3330 246256
rect 3386 246200 3391 246256
rect -960 246198 3391 246200
rect -960 246108 480 246198
rect 3325 246195 3391 246198
rect 499520 245836 500960 246076
rect -960 241484 480 241724
rect 499520 241484 500960 241724
rect 103421 238642 103487 238645
rect 103646 238642 103652 238644
rect 103376 238640 103652 238642
rect 103376 238584 103426 238640
rect 103482 238584 103652 238640
rect 103376 238582 103652 238584
rect 103421 238579 103487 238582
rect 103646 238580 103652 238582
rect 103716 238580 103722 238644
rect -960 237132 480 237372
rect 496261 237010 496327 237013
rect 499520 237010 500960 237100
rect 496261 237008 500960 237010
rect 496261 236952 496266 237008
rect 496322 236952 500960 237008
rect 496261 236950 500960 236952
rect 496261 236947 496327 236950
rect 499520 236860 500960 236950
rect 62481 236194 62547 236197
rect 62614 236194 62620 236196
rect 62481 236192 62620 236194
rect 62481 236136 62486 236192
rect 62542 236136 62620 236192
rect 62481 236134 62620 236136
rect 62481 236131 62547 236134
rect 62614 236132 62620 236134
rect 62684 236132 62690 236196
rect 61469 236060 61535 236061
rect 61469 236056 61516 236060
rect 61580 236058 61586 236060
rect 61469 236000 61474 236056
rect 61469 235996 61516 236000
rect 61580 235998 61626 236058
rect 61580 235996 61586 235998
rect 61469 235995 61535 235996
rect -960 232508 480 232748
rect 212390 232460 212396 232524
rect 212460 232522 212466 232524
rect 240317 232522 240383 232525
rect 212460 232520 240383 232522
rect 212460 232464 240322 232520
rect 240378 232464 240383 232520
rect 499520 232508 500960 232748
rect 212460 232462 240383 232464
rect 212460 232460 212466 232462
rect 240317 232459 240383 232462
rect 153469 229802 153535 229805
rect 188286 229802 188292 229804
rect 153469 229800 188292 229802
rect 153469 229744 153474 229800
rect 153530 229744 188292 229800
rect 153469 229742 188292 229744
rect 153469 229739 153535 229742
rect 188286 229740 188292 229742
rect 188356 229740 188362 229804
rect 103421 229124 103487 229125
rect 103421 229122 103468 229124
rect 103376 229120 103468 229122
rect 103532 229122 103538 229124
rect 103376 229064 103426 229120
rect 103376 229062 103468 229064
rect 103421 229060 103468 229062
rect 103532 229062 103614 229122
rect 103532 229060 103538 229062
rect 103421 229059 103487 229060
rect 103421 228988 103487 228989
rect 103421 228986 103468 228988
rect 103376 228984 103468 228986
rect 103532 228986 103538 228988
rect 103376 228928 103426 228984
rect 103376 228926 103468 228928
rect 103421 228924 103468 228926
rect 103532 228926 103614 228986
rect 103532 228924 103538 228926
rect 103421 228923 103487 228924
rect -960 228156 480 228396
rect 44030 228244 44036 228308
rect 44100 228306 44106 228308
rect 167453 228306 167519 228309
rect 44100 228304 167519 228306
rect 44100 228248 167458 228304
rect 167514 228248 167519 228304
rect 44100 228246 167519 228248
rect 44100 228244 44106 228246
rect 167453 228243 167519 228246
rect 53046 228108 53052 228172
rect 53116 228170 53122 228172
rect 167361 228170 167427 228173
rect 175825 228172 175891 228173
rect 175774 228170 175780 228172
rect 53116 228168 167427 228170
rect 53116 228112 167366 228168
rect 167422 228112 167427 228168
rect 53116 228110 167427 228112
rect 175734 228110 175780 228170
rect 175844 228168 175891 228172
rect 175886 228112 175891 228168
rect 53116 228108 53122 228110
rect 167361 228107 167427 228110
rect 175774 228108 175780 228110
rect 175844 228108 175891 228112
rect 175825 228107 175891 228108
rect 499520 227884 500960 228124
rect 135621 227084 135687 227085
rect 135621 227082 135668 227084
rect 135576 227080 135668 227082
rect 135732 227082 135738 227084
rect 136541 227082 136607 227085
rect 135732 227080 136607 227082
rect 135576 227024 135626 227080
rect 135732 227024 136546 227080
rect 136602 227024 136607 227080
rect 135576 227022 135668 227024
rect 135621 227020 135668 227022
rect 135732 227022 136607 227024
rect 135732 227020 135738 227022
rect 135621 227019 135687 227020
rect 136541 227019 136607 227022
rect 137185 226674 137251 226677
rect 138606 226674 138612 226676
rect 137185 226672 138612 226674
rect 137185 226616 137190 226672
rect 137246 226616 138612 226672
rect 137185 226614 138612 226616
rect 137185 226611 137251 226614
rect 138606 226612 138612 226614
rect 138676 226612 138682 226676
rect 103421 224908 103487 224909
rect 103421 224904 103468 224908
rect 103532 224906 103538 224908
rect 103421 224848 103426 224904
rect 103421 224844 103468 224848
rect 103532 224846 103578 224906
rect 103532 224844 103538 224846
rect 103421 224843 103487 224844
rect 63718 224436 63724 224500
rect 63788 224498 63794 224500
rect 100937 224498 101003 224501
rect 63788 224496 101003 224498
rect 63788 224440 100942 224496
rect 100998 224440 101003 224496
rect 63788 224438 101003 224440
rect 63788 224436 63794 224438
rect 100937 224435 101003 224438
rect -960 223954 480 224044
rect 3049 223954 3115 223957
rect -960 223952 3115 223954
rect -960 223896 3054 223952
rect 3110 223896 3115 223952
rect -960 223894 3115 223896
rect -960 223804 480 223894
rect 3049 223891 3115 223894
rect 289629 223684 289695 223685
rect 289629 223680 289676 223684
rect 289740 223682 289746 223684
rect 496537 223682 496603 223685
rect 499520 223682 500960 223772
rect 289629 223624 289634 223680
rect 289629 223620 289676 223624
rect 289740 223622 289786 223682
rect 496537 223680 500960 223682
rect 496537 223624 496542 223680
rect 496598 223624 500960 223680
rect 496537 223622 500960 223624
rect 289740 223620 289746 223622
rect 289629 223619 289695 223620
rect 496537 223619 496603 223622
rect 499520 223532 500960 223622
rect 255957 223274 256023 223277
rect 260741 223274 260807 223277
rect 255957 223272 260807 223274
rect 255957 223216 255962 223272
rect 256018 223216 260746 223272
rect 260802 223216 260807 223272
rect 255957 223214 260807 223216
rect 255957 223211 256023 223214
rect 260741 223211 260807 223214
rect 3325 222594 3391 222597
rect 240133 222594 240199 222597
rect 3325 222592 240199 222594
rect 3325 222536 3330 222592
rect 3386 222536 240138 222592
rect 240194 222536 240199 222592
rect 3325 222534 240199 222536
rect 3325 222531 3391 222534
rect 240133 222531 240199 222534
rect 214373 222458 214439 222461
rect 224718 222458 224724 222460
rect 214373 222456 224724 222458
rect 214373 222400 214378 222456
rect 214434 222400 224724 222456
rect 214373 222398 224724 222400
rect 214373 222395 214439 222398
rect 224718 222396 224724 222398
rect 224788 222396 224794 222460
rect 59118 222260 59124 222324
rect 59188 222322 59194 222324
rect 61837 222322 61903 222325
rect 59188 222320 61903 222322
rect 59188 222264 61842 222320
rect 61898 222264 61903 222320
rect 59188 222262 61903 222264
rect 59188 222260 59194 222262
rect 61837 222259 61903 222262
rect 75177 222322 75243 222325
rect 83958 222322 83964 222324
rect 75177 222320 83964 222322
rect 75177 222264 75182 222320
rect 75238 222264 83964 222320
rect 75177 222262 83964 222264
rect 75177 222259 75243 222262
rect 83958 222260 83964 222262
rect 84028 222260 84034 222324
rect 204110 222260 204116 222324
rect 204180 222322 204186 222324
rect 207381 222322 207447 222325
rect 204180 222320 207447 222322
rect 204180 222264 207386 222320
rect 207442 222264 207447 222320
rect 204180 222262 207447 222264
rect 204180 222260 204186 222262
rect 207381 222259 207447 222262
rect 209037 220828 209103 220829
rect 127566 220826 127572 220828
rect 122790 220766 127572 220826
rect 79317 220690 79383 220693
rect 122790 220690 122850 220766
rect 127566 220764 127572 220766
rect 127636 220764 127642 220828
rect 209037 220824 209084 220828
rect 209148 220826 209154 220828
rect 209037 220768 209042 220824
rect 209037 220764 209084 220768
rect 209148 220766 209194 220826
rect 209148 220764 209154 220766
rect 209037 220763 209103 220764
rect 79317 220688 122850 220690
rect 79317 220632 79322 220688
rect 79378 220632 122850 220688
rect 79317 220630 122850 220632
rect 123385 220690 123451 220693
rect 124806 220690 124812 220692
rect 123385 220688 124812 220690
rect 123385 220632 123390 220688
rect 123446 220632 124812 220688
rect 123385 220630 124812 220632
rect 79317 220627 79383 220630
rect 123385 220627 123451 220630
rect 124806 220628 124812 220630
rect 124876 220628 124882 220692
rect 259177 220690 259243 220693
rect 496169 220690 496235 220693
rect 259177 220688 496235 220690
rect 259177 220632 259182 220688
rect 259238 220632 496174 220688
rect 496230 220632 496235 220688
rect 259177 220630 496235 220632
rect 259177 220627 259243 220630
rect 496169 220627 496235 220630
rect 55029 220554 55095 220557
rect 373993 220554 374059 220557
rect 55029 220552 374059 220554
rect 55029 220496 55034 220552
rect 55090 220496 373998 220552
rect 374054 220496 374059 220552
rect 55029 220494 374059 220496
rect 55029 220491 55095 220494
rect 373993 220491 374059 220494
rect 213177 220420 213243 220421
rect 213126 220418 213132 220420
rect 213086 220358 213132 220418
rect 213196 220416 213243 220420
rect 213238 220360 213243 220416
rect 213126 220356 213132 220358
rect 213196 220356 213243 220360
rect 213177 220355 213243 220356
rect 159081 220282 159147 220285
rect 318241 220282 318307 220285
rect 159081 220280 318307 220282
rect 159081 220224 159086 220280
rect 159142 220224 318246 220280
rect 318302 220224 318307 220280
rect 159081 220222 318307 220224
rect 159081 220219 159147 220222
rect 318241 220219 318307 220222
rect 5441 220146 5507 220149
rect 311709 220146 311775 220149
rect 5441 220144 311775 220146
rect 5441 220088 5446 220144
rect 5502 220088 311714 220144
rect 311770 220088 311775 220144
rect 5441 220086 311775 220088
rect 5441 220083 5507 220086
rect 311709 220083 311775 220086
rect 34462 219948 34468 220012
rect 34532 220010 34538 220012
rect 34789 220010 34855 220013
rect 42057 220012 42123 220013
rect 42006 220010 42012 220012
rect 34532 220008 34855 220010
rect 34532 219952 34794 220008
rect 34850 219952 34855 220008
rect 34532 219950 34855 219952
rect 41966 219950 42012 220010
rect 42076 220008 42123 220012
rect 42118 219952 42123 220008
rect 34532 219948 34538 219950
rect 34789 219947 34855 219950
rect 42006 219948 42012 219950
rect 42076 219948 42123 219952
rect 42057 219947 42123 219948
rect 49969 220010 50035 220013
rect 51574 220010 51580 220012
rect 49969 220008 51580 220010
rect 49969 219952 49974 220008
rect 50030 219952 51580 220008
rect 49969 219950 51580 219952
rect 49969 219947 50035 219950
rect 51574 219948 51580 219950
rect 51644 219948 51650 220012
rect 54334 219948 54340 220012
rect 54404 220010 54410 220012
rect 54661 220010 54727 220013
rect 54404 220008 54727 220010
rect 54404 219952 54666 220008
rect 54722 219952 54727 220008
rect 54404 219950 54727 219952
rect 54404 219948 54410 219950
rect 54661 219947 54727 219950
rect 68134 219948 68140 220012
rect 68204 220010 68210 220012
rect 68277 220010 68343 220013
rect 68204 220008 68343 220010
rect 68204 219952 68282 220008
rect 68338 219952 68343 220008
rect 68204 219950 68343 219952
rect 68204 219948 68210 219950
rect 68277 219947 68343 219950
rect 79409 220010 79475 220013
rect 94497 220012 94563 220013
rect 79542 220010 79548 220012
rect 79409 220008 79548 220010
rect 79409 219952 79414 220008
rect 79470 219952 79548 220008
rect 79409 219950 79548 219952
rect 79409 219947 79475 219950
rect 79542 219948 79548 219950
rect 79612 219948 79618 220012
rect 94446 220010 94452 220012
rect 94406 219950 94452 220010
rect 94516 220008 94563 220012
rect 94558 219952 94563 220008
rect 94446 219948 94452 219950
rect 94516 219948 94563 219952
rect 101254 219948 101260 220012
rect 101324 220010 101330 220012
rect 101397 220010 101463 220013
rect 101324 220008 101463 220010
rect 101324 219952 101402 220008
rect 101458 219952 101463 220008
rect 101324 219950 101463 219952
rect 101324 219948 101330 219950
rect 94497 219947 94563 219948
rect 101397 219947 101463 219950
rect 134374 219948 134380 220012
rect 134444 220010 134450 220012
rect 134517 220010 134583 220013
rect 134444 220008 134583 220010
rect 134444 219952 134522 220008
rect 134578 219952 134583 220008
rect 134444 219950 134583 219952
rect 134444 219948 134450 219950
rect 134517 219947 134583 219950
rect 153694 219948 153700 220012
rect 153764 220010 153770 220012
rect 154021 220010 154087 220013
rect 153764 220008 154087 220010
rect 153764 219952 154026 220008
rect 154082 219952 154087 220008
rect 153764 219950 154087 219952
rect 153764 219948 153770 219950
rect 154021 219947 154087 219950
rect 186814 219948 186820 220012
rect 186884 220010 186890 220012
rect 187141 220010 187207 220013
rect 186884 220008 187207 220010
rect 186884 219952 187146 220008
rect 187202 219952 187207 220008
rect 186884 219950 187207 219952
rect 186884 219948 186890 219950
rect 187141 219947 187207 219950
rect 193070 219948 193076 220012
rect 193140 220010 193146 220012
rect 193765 220010 193831 220013
rect 226977 220012 227043 220013
rect 226926 220010 226932 220012
rect 193140 220008 193831 220010
rect 193140 219952 193770 220008
rect 193826 219952 193831 220008
rect 193140 219950 193831 219952
rect 226886 219950 226932 220010
rect 226996 220008 227043 220012
rect 227038 219952 227043 220008
rect 193140 219948 193146 219950
rect 193765 219947 193831 219950
rect 226926 219948 226932 219950
rect 226996 219948 227043 219952
rect 226977 219947 227043 219948
rect 235257 220010 235323 220013
rect 243486 220010 243492 220012
rect 235257 220008 243492 220010
rect 235257 219952 235262 220008
rect 235318 219952 243492 220008
rect 235257 219950 243492 219952
rect 235257 219947 235323 219950
rect 243486 219948 243492 219950
rect 243556 219948 243562 220012
rect 253054 219948 253060 220012
rect 253124 220010 253130 220012
rect 253381 220010 253447 220013
rect 253124 220008 253447 220010
rect 253124 219952 253386 220008
rect 253442 219952 253447 220008
rect 253124 219950 253447 219952
rect 253124 219948 253130 219950
rect 253381 219947 253447 219950
rect 280521 220010 280587 220013
rect 280654 220010 280660 220012
rect 280521 220008 280660 220010
rect 280521 219952 280526 220008
rect 280582 219952 280660 220008
rect 280521 219950 280660 219952
rect 280521 219947 280587 219950
rect 280654 219948 280660 219950
rect 280724 219948 280730 220012
rect 77886 219812 77892 219876
rect 77956 219874 77962 219876
rect 257705 219874 257771 219877
rect 77956 219872 257771 219874
rect 77956 219816 257710 219872
rect 257766 219816 257771 219872
rect 77956 219814 257771 219816
rect 77956 219812 77962 219814
rect 257705 219811 257771 219814
rect 264973 219874 265039 219877
rect 266629 219874 266695 219877
rect 264973 219872 266695 219874
rect 264973 219816 264978 219872
rect 265034 219816 266634 219872
rect 266690 219816 266695 219872
rect 264973 219814 266695 219816
rect 264973 219811 265039 219814
rect 266629 219811 266695 219814
rect 77753 219738 77819 219741
rect 240133 219740 240199 219741
rect 80646 219738 80652 219740
rect 77753 219736 80652 219738
rect 77753 219680 77758 219736
rect 77814 219680 80652 219736
rect 77753 219678 80652 219680
rect 77753 219675 77819 219678
rect 80646 219676 80652 219678
rect 80716 219676 80722 219740
rect 240133 219736 240180 219740
rect 240244 219738 240250 219740
rect 240133 219680 240138 219736
rect 240133 219676 240180 219680
rect 240244 219678 240290 219738
rect 240244 219676 240250 219678
rect 240133 219675 240199 219676
rect 162526 219540 162532 219604
rect 162596 219602 162602 219604
rect 162761 219602 162827 219605
rect 162596 219600 162827 219602
rect 162596 219544 162766 219600
rect 162822 219544 162827 219600
rect 162596 219542 162827 219544
rect 162596 219540 162602 219542
rect 162761 219539 162827 219542
rect 205030 219540 205036 219604
rect 205100 219602 205106 219604
rect 205173 219602 205239 219605
rect 205100 219600 205239 219602
rect 205100 219544 205178 219600
rect 205234 219544 205239 219600
rect 205100 219542 205239 219544
rect 205100 219540 205106 219542
rect 205173 219539 205239 219542
rect -960 219330 480 219420
rect 87454 219404 87460 219468
rect 87524 219466 87530 219468
rect 87781 219466 87847 219469
rect 87524 219464 87847 219466
rect 87524 219408 87786 219464
rect 87842 219408 87847 219464
rect 87524 219406 87847 219408
rect 87524 219404 87530 219406
rect 87781 219403 87847 219406
rect 96613 219468 96679 219469
rect 96613 219464 96660 219468
rect 96724 219466 96730 219468
rect 114921 219466 114987 219469
rect 115054 219466 115060 219468
rect 96613 219408 96618 219464
rect 96613 219404 96660 219408
rect 96724 219406 96770 219466
rect 114921 219464 115060 219466
rect 114921 219408 114926 219464
rect 114982 219408 115060 219464
rect 114921 219406 115060 219408
rect 96724 219404 96730 219406
rect 96613 219403 96679 219404
rect 114921 219403 114987 219406
rect 115054 219404 115060 219406
rect 115124 219404 115130 219468
rect 161289 219466 161355 219469
rect 162894 219466 162900 219468
rect 161289 219464 162900 219466
rect 161289 219408 161294 219464
rect 161350 219408 162900 219464
rect 161289 219406 162900 219408
rect 161289 219403 161355 219406
rect 162894 219404 162900 219406
rect 162964 219404 162970 219468
rect 167913 219466 167979 219469
rect 173985 219468 174051 219469
rect 172462 219466 172468 219468
rect 167913 219464 172468 219466
rect 167913 219408 167918 219464
rect 167974 219408 172468 219464
rect 167913 219406 172468 219408
rect 167913 219403 167979 219406
rect 172462 219404 172468 219406
rect 172532 219404 172538 219468
rect 173934 219466 173940 219468
rect 173894 219406 173940 219466
rect 174004 219464 174051 219468
rect 174046 219408 174051 219464
rect 173934 219404 173940 219406
rect 174004 219404 174051 219408
rect 173985 219403 174051 219404
rect 181161 219466 181227 219469
rect 184974 219466 184980 219468
rect 181161 219464 184980 219466
rect 181161 219408 181166 219464
rect 181222 219408 184980 219464
rect 181161 219406 184980 219408
rect 181161 219403 181227 219406
rect 184974 219404 184980 219406
rect 185044 219404 185050 219468
rect 234153 219466 234219 219469
rect 235942 219466 235948 219468
rect 234153 219464 235948 219466
rect 234153 219408 234158 219464
rect 234214 219408 235948 219464
rect 234153 219406 235948 219408
rect 234153 219403 234219 219406
rect 235942 219404 235948 219406
rect 236012 219404 236018 219468
rect 273110 219404 273116 219468
rect 273180 219466 273186 219468
rect 273253 219466 273319 219469
rect 293217 219468 293283 219469
rect 293166 219466 293172 219468
rect 273180 219464 273319 219466
rect 273180 219408 273258 219464
rect 273314 219408 273319 219464
rect 273180 219406 273319 219408
rect 293126 219406 293172 219466
rect 293236 219464 293283 219468
rect 293278 219408 293283 219464
rect 273180 219404 273186 219406
rect 273253 219403 273319 219406
rect 293166 219404 293172 219406
rect 293236 219404 293283 219408
rect 293217 219403 293283 219404
rect 3601 219330 3667 219333
rect -960 219328 3667 219330
rect -960 219272 3606 219328
rect 3662 219272 3667 219328
rect -960 219270 3667 219272
rect -960 219180 480 219270
rect 3601 219267 3667 219270
rect 219382 219268 219388 219332
rect 219452 219330 219458 219332
rect 220261 219330 220327 219333
rect 244917 219330 244983 219333
rect 219452 219328 220327 219330
rect 219452 219272 220266 219328
rect 220322 219272 220327 219328
rect 219452 219270 220327 219272
rect 219452 219268 219458 219270
rect 220261 219267 220327 219270
rect 238710 219328 244983 219330
rect 238710 219272 244922 219328
rect 244978 219272 244983 219328
rect 238710 219270 244983 219272
rect 209998 218588 210004 218652
rect 210068 218650 210074 218652
rect 238710 218650 238770 219270
rect 244917 219267 244983 219270
rect 495433 219058 495499 219061
rect 499520 219058 500960 219148
rect 495433 219056 500960 219058
rect 495433 219000 495438 219056
rect 495494 219000 500960 219056
rect 495433 218998 500960 219000
rect 495433 218995 495499 218998
rect 499520 218908 500960 218998
rect 210068 218590 238770 218650
rect 210068 218588 210074 218590
rect 9489 217834 9555 217837
rect 10182 217834 10242 217940
rect 9489 217832 10242 217834
rect 9489 217776 9494 217832
rect 9550 217776 10242 217832
rect 9489 217774 10242 217776
rect 9489 217771 9555 217774
rect -960 214978 480 215068
rect 3601 214978 3667 214981
rect 312445 214978 312511 214981
rect 312629 214978 312695 214981
rect -960 214976 3667 214978
rect -960 214920 3606 214976
rect 3662 214920 3667 214976
rect -960 214918 3667 214920
rect 309948 214976 312695 214978
rect 309948 214920 312450 214976
rect 312506 214920 312634 214976
rect 312690 214920 312695 214976
rect 309948 214918 312695 214920
rect -960 214828 480 214918
rect 3601 214915 3667 214918
rect 312445 214915 312511 214918
rect 312629 214915 312695 214918
rect 499520 214556 500960 214796
rect -960 210204 480 210444
rect 499520 209932 500960 210172
rect 8017 208314 8083 208317
rect 8017 208312 10058 208314
rect 8017 208256 8022 208312
rect 8078 208256 10058 208312
rect 8017 208254 10058 208256
rect 8017 208251 8083 208254
rect 9998 208148 10058 208254
rect -960 206002 480 206092
rect 2865 206002 2931 206005
rect -960 206000 2931 206002
rect -960 205944 2870 206000
rect 2926 205944 2931 206000
rect -960 205942 2931 205944
rect -960 205852 480 205942
rect 2865 205939 2931 205942
rect 496169 205730 496235 205733
rect 499520 205730 500960 205820
rect 496169 205728 500960 205730
rect 496169 205672 496174 205728
rect 496230 205672 500960 205728
rect 496169 205670 500960 205672
rect 496169 205667 496235 205670
rect 499520 205580 500960 205670
rect 312077 205186 312143 205189
rect 312537 205186 312603 205189
rect 309948 205184 312603 205186
rect 309948 205128 312082 205184
rect 312138 205128 312542 205184
rect 312598 205128 312603 205184
rect 309948 205126 312603 205128
rect 312077 205123 312143 205126
rect 312537 205123 312603 205126
rect -960 201378 480 201468
rect 3233 201378 3299 201381
rect -960 201376 3299 201378
rect -960 201320 3238 201376
rect 3294 201320 3299 201376
rect -960 201318 3299 201320
rect -960 201228 480 201318
rect 3233 201315 3299 201318
rect 495433 201106 495499 201109
rect 499520 201106 500960 201196
rect 495433 201104 500960 201106
rect 495433 201048 495438 201104
rect 495494 201048 500960 201104
rect 495433 201046 500960 201048
rect 495433 201043 495499 201046
rect 499520 200956 500960 201046
rect 7373 197842 7439 197845
rect 10182 197842 10242 198356
rect 7373 197840 10242 197842
rect 7373 197784 7378 197840
rect 7434 197784 10242 197840
rect 7373 197782 10242 197784
rect 7373 197779 7439 197782
rect -960 196876 480 197116
rect 495433 196754 495499 196757
rect 499520 196754 500960 196844
rect 495433 196752 500960 196754
rect 495433 196696 495438 196752
rect 495494 196696 500960 196752
rect 495433 196694 500960 196696
rect 495433 196691 495499 196694
rect 499520 196604 500960 196694
rect 312905 195394 312971 195397
rect 309948 195392 312971 195394
rect 309948 195336 312910 195392
rect 312966 195336 312971 195392
rect 309948 195334 312971 195336
rect 312905 195331 312971 195334
rect -960 192252 480 192492
rect 495433 192130 495499 192133
rect 499520 192130 500960 192220
rect 495433 192128 500960 192130
rect 495433 192072 495438 192128
rect 495494 192072 500960 192128
rect 495433 192070 500960 192072
rect 495433 192067 495499 192070
rect 499520 191980 500960 192070
rect 8201 189002 8267 189005
rect 8201 189000 10058 189002
rect 8201 188944 8206 189000
rect 8262 188944 10058 189000
rect 8201 188942 10058 188944
rect 8201 188939 8267 188942
rect 9998 188564 10058 188942
rect -960 188050 480 188140
rect 3325 188050 3391 188053
rect -960 188048 3391 188050
rect -960 187992 3330 188048
rect 3386 187992 3391 188048
rect -960 187990 3391 187992
rect -960 187900 480 187990
rect 3325 187987 3391 187990
rect 495433 187778 495499 187781
rect 499520 187778 500960 187868
rect 495433 187776 500960 187778
rect 495433 187720 495438 187776
rect 495494 187720 500960 187776
rect 495433 187718 500960 187720
rect 495433 187715 495499 187718
rect 499520 187628 500960 187718
rect 312169 185602 312235 185605
rect 312445 185602 312511 185605
rect 309948 185600 312511 185602
rect 309948 185544 312174 185600
rect 312230 185544 312450 185600
rect 312506 185544 312511 185600
rect 309948 185542 312511 185544
rect 312169 185539 312235 185542
rect 312445 185539 312511 185542
rect -960 183426 480 183516
rect 3049 183426 3115 183429
rect -960 183424 3115 183426
rect -960 183368 3054 183424
rect 3110 183368 3115 183424
rect -960 183366 3115 183368
rect -960 183276 480 183366
rect 3049 183363 3115 183366
rect 496353 183426 496419 183429
rect 499520 183426 500960 183516
rect 496353 183424 500960 183426
rect 496353 183368 496358 183424
rect 496414 183368 500960 183424
rect 496353 183366 500960 183368
rect 496353 183363 496419 183366
rect 499520 183276 500960 183366
rect -960 179074 480 179164
rect 3325 179074 3391 179077
rect -960 179072 3391 179074
rect -960 179016 3330 179072
rect 3386 179016 3391 179072
rect -960 179014 3391 179016
rect -960 178924 480 179014
rect 3325 179011 3391 179014
rect 7465 178938 7531 178941
rect 7465 178936 10058 178938
rect 7465 178880 7470 178936
rect 7526 178880 10058 178936
rect 7465 178878 10058 178880
rect 7465 178875 7531 178878
rect 9998 178772 10058 178878
rect 496629 178802 496695 178805
rect 499520 178802 500960 178892
rect 496629 178800 500960 178802
rect 496629 178744 496634 178800
rect 496690 178744 500960 178800
rect 496629 178742 500960 178744
rect 496629 178739 496695 178742
rect 499520 178652 500960 178742
rect 312353 175810 312419 175813
rect 309948 175808 312419 175810
rect 309948 175752 312358 175808
rect 312414 175752 312419 175808
rect 309948 175750 312419 175752
rect 312353 175747 312419 175750
rect -960 174300 480 174540
rect 495433 174450 495499 174453
rect 499520 174450 500960 174540
rect 495433 174448 500960 174450
rect 495433 174392 495438 174448
rect 495494 174392 500960 174448
rect 495433 174390 500960 174392
rect 495433 174387 495499 174390
rect 499520 174300 500960 174390
rect -960 169948 480 170188
rect 496721 169826 496787 169829
rect 499520 169826 500960 169916
rect 496721 169824 500960 169826
rect 496721 169768 496726 169824
rect 496782 169768 500960 169824
rect 496721 169766 500960 169768
rect 496721 169763 496787 169766
rect 499520 169676 500960 169766
rect 7373 168466 7439 168469
rect 10182 168466 10242 168980
rect 7373 168464 10242 168466
rect 7373 168408 7378 168464
rect 7434 168408 10242 168464
rect 7373 168406 10242 168408
rect 7373 168403 7439 168406
rect 312077 166018 312143 166021
rect 309948 166016 312143 166018
rect 309948 165960 312082 166016
rect 312138 165960 312143 166016
rect 309948 165958 312143 165960
rect 312077 165955 312143 165958
rect -960 165596 480 165836
rect 499520 165324 500960 165564
rect -960 161122 480 161212
rect 3325 161122 3391 161125
rect -960 161120 3391 161122
rect -960 161064 3330 161120
rect 3386 161064 3391 161120
rect -960 161062 3391 161064
rect -960 160972 480 161062
rect 3325 161059 3391 161062
rect 499520 160700 500960 160940
rect 7005 158810 7071 158813
rect 10182 158810 10242 159188
rect 7005 158808 10242 158810
rect 7005 158752 7010 158808
rect 7066 158752 10242 158808
rect 7005 158750 10242 158752
rect 7005 158747 7071 158750
rect -960 156770 480 156860
rect 3141 156770 3207 156773
rect -960 156768 3207 156770
rect -960 156712 3146 156768
rect 3202 156712 3207 156768
rect -960 156710 3207 156712
rect -960 156620 480 156710
rect 3141 156707 3207 156710
rect 499520 156348 500960 156588
rect 312169 156226 312235 156229
rect 309948 156224 312235 156226
rect 309948 156168 312174 156224
rect 312230 156168 312235 156224
rect 309948 156166 312235 156168
rect 312169 156163 312235 156166
rect -960 152146 480 152236
rect 4061 152146 4127 152149
rect -960 152144 4127 152146
rect -960 152088 4066 152144
rect 4122 152088 4127 152144
rect -960 152086 4127 152088
rect -960 151996 480 152086
rect 4061 152083 4127 152086
rect 499520 151724 500960 151964
rect 6913 149154 6979 149157
rect 7557 149154 7623 149157
rect 10182 149154 10242 149396
rect 6913 149152 10242 149154
rect 6913 149096 6918 149152
rect 6974 149096 7562 149152
rect 7618 149096 10242 149152
rect 6913 149094 10242 149096
rect 6913 149091 6979 149094
rect 7557 149091 7623 149094
rect -960 147644 480 147884
rect 495525 147522 495591 147525
rect 499520 147522 500960 147612
rect 495525 147520 500960 147522
rect 495525 147464 495530 147520
rect 495586 147464 500960 147520
rect 495525 147462 500960 147464
rect 495525 147459 495591 147462
rect 499520 147372 500960 147462
rect 312261 146434 312327 146437
rect 312721 146434 312787 146437
rect 309948 146432 312787 146434
rect 309948 146376 312266 146432
rect 312322 146376 312726 146432
rect 312782 146376 312787 146432
rect 309948 146374 312787 146376
rect 312261 146371 312327 146374
rect 312721 146371 312787 146374
rect -960 143170 480 143260
rect 3969 143170 4035 143173
rect -960 143168 4035 143170
rect -960 143112 3974 143168
rect 4030 143112 4035 143168
rect -960 143110 4035 143112
rect -960 143020 480 143110
rect 3969 143107 4035 143110
rect 495433 142898 495499 142901
rect 499520 142898 500960 142988
rect 495433 142896 500960 142898
rect 495433 142840 495438 142896
rect 495494 142840 500960 142896
rect 495433 142838 500960 142840
rect 495433 142835 495499 142838
rect 499520 142748 500960 142838
rect 7649 139770 7715 139773
rect 7649 139768 10058 139770
rect 7649 139712 7654 139768
rect 7710 139712 10058 139768
rect 7649 139710 10058 139712
rect 7649 139707 7715 139710
rect 9998 139604 10058 139710
rect -960 138818 480 138908
rect 3325 138818 3391 138821
rect -960 138816 3391 138818
rect -960 138760 3330 138816
rect 3386 138760 3391 138816
rect -960 138758 3391 138760
rect -960 138668 480 138758
rect 3325 138755 3391 138758
rect 499520 138396 500960 138636
rect 312813 136642 312879 136645
rect 309948 136640 312879 136642
rect 309948 136584 312818 136640
rect 312874 136584 312879 136640
rect 309948 136582 312879 136584
rect 312813 136579 312879 136582
rect -960 134194 480 134284
rect 4061 134194 4127 134197
rect -960 134192 4127 134194
rect -960 134136 4066 134192
rect 4122 134136 4127 134192
rect -960 134134 4127 134136
rect -960 134044 480 134134
rect 4061 134131 4127 134134
rect 499520 133772 500960 134012
rect 8201 129978 8267 129981
rect 8201 129976 10058 129978
rect -960 129842 480 129932
rect 8201 129920 8206 129976
rect 8262 129920 10058 129976
rect 8201 129918 10058 129920
rect 8201 129915 8267 129918
rect 4061 129842 4127 129845
rect -960 129840 4127 129842
rect -960 129784 4066 129840
rect 4122 129784 4127 129840
rect 9998 129812 10058 129918
rect -960 129782 4127 129784
rect -960 129692 480 129782
rect 4061 129779 4127 129782
rect 496353 129570 496419 129573
rect 499520 129570 500960 129660
rect 496353 129568 500960 129570
rect 496353 129512 496358 129568
rect 496414 129512 500960 129568
rect 496353 129510 500960 129512
rect 496353 129507 496419 129510
rect 499520 129420 500960 129510
rect 312261 126850 312327 126853
rect 309948 126848 312327 126850
rect 309948 126792 312266 126848
rect 312322 126792 312327 126848
rect 309948 126790 312327 126792
rect 312261 126787 312327 126790
rect -960 125218 480 125308
rect 3969 125218 4035 125221
rect -960 125216 4035 125218
rect -960 125160 3974 125216
rect 4030 125160 4035 125216
rect -960 125158 4035 125160
rect -960 125068 480 125158
rect 3969 125155 4035 125158
rect 499520 125068 500960 125308
rect 8937 121410 9003 121413
rect 219014 121410 219020 121412
rect 8937 121408 219020 121410
rect 8937 121352 8942 121408
rect 8998 121352 219020 121408
rect 8937 121350 219020 121352
rect 8937 121347 9003 121350
rect 219014 121348 219020 121350
rect 219084 121410 219090 121412
rect 219566 121410 219572 121412
rect 219084 121350 219572 121410
rect 219084 121348 219090 121350
rect 219566 121348 219572 121350
rect 219636 121348 219642 121412
rect -960 120866 480 120956
rect 2773 120866 2839 120869
rect -960 120864 2839 120866
rect -960 120808 2778 120864
rect 2834 120808 2839 120864
rect -960 120806 2839 120808
rect -960 120716 480 120806
rect 2773 120803 2839 120806
rect 43529 120730 43595 120733
rect 96429 120732 96495 120733
rect 44030 120730 44036 120732
rect 43529 120728 44036 120730
rect 43529 120672 43534 120728
rect 43590 120672 44036 120728
rect 43529 120670 44036 120672
rect 43529 120667 43595 120670
rect 44030 120668 44036 120670
rect 44100 120668 44106 120732
rect 96429 120730 96476 120732
rect 96384 120728 96476 120730
rect 96384 120672 96434 120728
rect 96384 120670 96476 120672
rect 96429 120668 96476 120670
rect 96540 120668 96546 120732
rect 103145 120730 103211 120733
rect 103278 120730 103284 120732
rect 103145 120728 103284 120730
rect 103145 120672 103150 120728
rect 103206 120672 103284 120728
rect 103145 120670 103284 120672
rect 96429 120667 96495 120668
rect 103145 120667 103211 120670
rect 103278 120668 103284 120670
rect 103348 120668 103354 120732
rect 116393 120730 116459 120733
rect 117078 120730 117084 120732
rect 116393 120728 117084 120730
rect 116393 120672 116398 120728
rect 116454 120672 117084 120728
rect 116393 120670 117084 120672
rect 116393 120667 116459 120670
rect 117078 120668 117084 120670
rect 117148 120668 117154 120732
rect 499520 120444 500960 120684
rect 34278 119988 34284 120052
rect 34348 120050 34354 120052
rect 34973 120050 35039 120053
rect 34348 120048 35039 120050
rect 34348 119992 34978 120048
rect 35034 119992 35039 120048
rect 34348 119990 35039 119992
rect 34348 119988 34354 119990
rect 34973 119987 35039 119990
rect 38745 120050 38811 120053
rect 38878 120050 38884 120052
rect 38745 120048 38884 120050
rect 38745 119992 38750 120048
rect 38806 119992 38884 120048
rect 38745 119990 38884 119992
rect 38745 119987 38811 119990
rect 38878 119988 38884 119990
rect 38948 119988 38954 120052
rect 55438 119988 55444 120052
rect 55508 120050 55514 120052
rect 63493 120050 63559 120053
rect 55508 120048 63559 120050
rect 55508 119992 63498 120048
rect 63554 119992 63559 120048
rect 55508 119990 63559 119992
rect 55508 119988 55514 119990
rect 63493 119987 63559 119990
rect 63677 120052 63743 120053
rect 63677 120048 63724 120052
rect 63788 120050 63794 120052
rect 63677 119992 63682 120048
rect 63677 119988 63724 119992
rect 63788 119990 63834 120050
rect 63788 119988 63794 119990
rect 131614 119988 131620 120052
rect 131684 120050 131690 120052
rect 161013 120050 161079 120053
rect 131684 120048 161079 120050
rect 131684 119992 161018 120048
rect 161074 119992 161079 120048
rect 131684 119990 161079 119992
rect 131684 119988 131690 119990
rect 63677 119987 63743 119988
rect 161013 119987 161079 119990
rect 172697 120050 172763 120053
rect 258022 120050 258028 120052
rect 172697 120048 258028 120050
rect 172697 119992 172702 120048
rect 172758 119992 258028 120048
rect 172697 119990 258028 119992
rect 172697 119987 172763 119990
rect 258022 119988 258028 119990
rect 258092 119988 258098 120052
rect 35157 119914 35223 119917
rect 162485 119916 162551 119917
rect 143206 119914 143212 119916
rect 35157 119912 143212 119914
rect 35157 119856 35162 119912
rect 35218 119856 143212 119912
rect 35157 119854 143212 119856
rect 35157 119851 35223 119854
rect 143206 119852 143212 119854
rect 143276 119852 143282 119916
rect 162485 119912 162532 119916
rect 162596 119914 162602 119916
rect 162485 119856 162490 119912
rect 162485 119852 162532 119856
rect 162596 119854 162642 119914
rect 162596 119852 162602 119854
rect 200614 119852 200620 119916
rect 200684 119914 200690 119916
rect 290457 119914 290523 119917
rect 200684 119912 290523 119914
rect 200684 119856 290462 119912
rect 290518 119856 290523 119912
rect 200684 119854 290523 119856
rect 200684 119852 200690 119854
rect 162485 119851 162551 119852
rect 290457 119851 290523 119854
rect 62614 119716 62620 119780
rect 62684 119778 62690 119780
rect 215753 119778 215819 119781
rect 62684 119776 215819 119778
rect 62684 119720 215758 119776
rect 215814 119720 215819 119776
rect 62684 119718 215819 119720
rect 62684 119716 62690 119718
rect 215753 119715 215819 119718
rect 61510 119580 61516 119644
rect 61580 119642 61586 119644
rect 215569 119642 215635 119645
rect 219198 119642 219204 119644
rect 61580 119640 215635 119642
rect 61580 119584 215574 119640
rect 215630 119584 215635 119640
rect 61580 119582 215635 119584
rect 61580 119580 61586 119582
rect 215569 119579 215635 119582
rect 215710 119582 219204 119642
rect 35341 119506 35407 119509
rect 215710 119506 215770 119582
rect 219198 119580 219204 119582
rect 219268 119580 219274 119644
rect 253933 119642 253999 119645
rect 254485 119642 254551 119645
rect 253933 119640 254551 119642
rect 253933 119584 253938 119640
rect 253994 119584 254490 119640
rect 254546 119584 254551 119640
rect 253933 119582 254551 119584
rect 253933 119579 253999 119582
rect 254485 119579 254551 119582
rect 216029 119508 216095 119509
rect 216029 119506 216076 119508
rect 35341 119504 215770 119506
rect 35341 119448 35346 119504
rect 35402 119448 215770 119504
rect 35341 119446 215770 119448
rect 215984 119504 216076 119506
rect 215984 119448 216034 119504
rect 215984 119446 216076 119448
rect 35341 119443 35407 119446
rect 216029 119444 216076 119446
rect 216140 119444 216146 119508
rect 289721 119506 289787 119509
rect 292113 119506 292179 119509
rect 289721 119504 292179 119506
rect 289721 119448 289726 119504
rect 289782 119448 292118 119504
rect 292174 119448 292179 119504
rect 289721 119446 292179 119448
rect 216029 119443 216095 119444
rect 289721 119443 289787 119446
rect 292113 119443 292179 119446
rect 34881 119370 34947 119373
rect 40534 119370 40540 119372
rect 34881 119368 40540 119370
rect 34881 119312 34886 119368
rect 34942 119312 40540 119368
rect 34881 119310 40540 119312
rect 34881 119307 34947 119310
rect 40534 119308 40540 119310
rect 40604 119308 40610 119372
rect 64045 119370 64111 119373
rect 228582 119370 228588 119372
rect 64045 119368 228588 119370
rect 64045 119312 64050 119368
rect 64106 119312 228588 119368
rect 64045 119310 228588 119312
rect 64045 119307 64111 119310
rect 228582 119308 228588 119310
rect 228652 119308 228658 119372
rect 254209 119370 254275 119373
rect 263726 119370 263732 119372
rect 254209 119368 263732 119370
rect 254209 119312 254214 119368
rect 254270 119312 263732 119368
rect 254209 119310 263732 119312
rect 254209 119307 254275 119310
rect 263726 119308 263732 119310
rect 263796 119308 263802 119372
rect 48129 119236 48195 119237
rect 48078 119234 48084 119236
rect 48038 119174 48084 119234
rect 48148 119232 48195 119236
rect 48190 119176 48195 119232
rect 48078 119172 48084 119174
rect 48148 119172 48195 119176
rect 104014 119172 104020 119236
rect 104084 119234 104090 119236
rect 238753 119234 238819 119237
rect 104084 119232 238819 119234
rect 104084 119176 238758 119232
rect 238814 119176 238819 119232
rect 104084 119174 238819 119176
rect 104084 119172 104090 119174
rect 48129 119171 48195 119172
rect 238753 119171 238819 119174
rect 34605 119098 34671 119101
rect 36486 119098 36492 119100
rect 34605 119096 36492 119098
rect 34605 119040 34610 119096
rect 34666 119040 36492 119096
rect 34605 119038 36492 119040
rect 34605 119035 34671 119038
rect 36486 119036 36492 119038
rect 36556 119036 36562 119100
rect 38837 119098 38903 119101
rect 135662 119098 135668 119100
rect 38837 119096 135668 119098
rect 38837 119040 38842 119096
rect 38898 119040 135668 119096
rect 38837 119038 135668 119040
rect 38837 119035 38903 119038
rect 135662 119036 135668 119038
rect 135732 119036 135738 119100
rect 145649 119098 145715 119101
rect 157517 119100 157583 119101
rect 215845 119100 215911 119101
rect 145782 119098 145788 119100
rect 145649 119096 145788 119098
rect 145649 119040 145654 119096
rect 145710 119040 145788 119096
rect 145649 119038 145788 119040
rect 145649 119035 145715 119038
rect 145782 119036 145788 119038
rect 145852 119036 145858 119100
rect 157517 119096 157564 119100
rect 157628 119098 157634 119100
rect 215845 119098 215892 119100
rect 157517 119040 157522 119096
rect 157517 119036 157564 119040
rect 157628 119038 157674 119098
rect 215800 119096 215892 119098
rect 215956 119098 215962 119100
rect 216581 119098 216647 119101
rect 215956 119096 216647 119098
rect 215800 119040 215850 119096
rect 215956 119040 216586 119096
rect 216642 119040 216647 119096
rect 215800 119038 215892 119040
rect 157628 119036 157634 119038
rect 215845 119036 215892 119038
rect 215956 119038 216647 119040
rect 215956 119036 215962 119038
rect 157517 119035 157583 119036
rect 215845 119035 215911 119036
rect 216581 119035 216647 119038
rect 34789 118962 34855 118965
rect 282678 118962 282684 118964
rect 34789 118960 282684 118962
rect 34789 118904 34794 118960
rect 34850 118904 282684 118960
rect 34789 118902 282684 118904
rect 34789 118899 34855 118902
rect 282678 118900 282684 118902
rect 282748 118900 282754 118964
rect 34881 118826 34947 118829
rect 35014 118826 35020 118828
rect 34881 118824 35020 118826
rect 34881 118768 34886 118824
rect 34942 118768 35020 118824
rect 34881 118766 35020 118768
rect 34881 118763 34947 118766
rect 35014 118764 35020 118766
rect 35084 118826 35090 118828
rect 48814 118826 48820 118828
rect 35084 118766 48820 118826
rect 35084 118764 35090 118766
rect 48814 118764 48820 118766
rect 48884 118764 48890 118828
rect 145741 118826 145807 118829
rect 147070 118826 147076 118828
rect 145741 118824 147076 118826
rect 145741 118768 145746 118824
rect 145802 118768 147076 118824
rect 145741 118766 147076 118768
rect 145741 118763 145807 118766
rect 147070 118764 147076 118766
rect 147140 118764 147146 118828
rect 261334 118628 261340 118692
rect 261404 118690 261410 118692
rect 261477 118690 261543 118693
rect 261404 118688 261543 118690
rect 261404 118632 261482 118688
rect 261538 118632 261543 118688
rect 261404 118630 261543 118632
rect 261404 118628 261410 118630
rect 261477 118627 261543 118630
rect 49877 118554 49943 118557
rect 234654 118554 234660 118556
rect 49877 118552 234660 118554
rect 49877 118496 49882 118552
rect 49938 118496 234660 118552
rect 49877 118494 234660 118496
rect 49877 118491 49943 118494
rect 234654 118492 234660 118494
rect 234724 118492 234730 118556
rect 235625 118554 235691 118557
rect 295374 118554 295380 118556
rect 235625 118552 295380 118554
rect 235625 118496 235630 118552
rect 235686 118496 295380 118552
rect 235625 118494 295380 118496
rect 235625 118491 235691 118494
rect 295374 118492 295380 118494
rect 295444 118492 295450 118556
rect 32438 118356 32444 118420
rect 32508 118418 32514 118420
rect 109125 118418 109191 118421
rect 32508 118416 109191 118418
rect 32508 118360 109130 118416
rect 109186 118360 109191 118416
rect 32508 118358 109191 118360
rect 32508 118356 32514 118358
rect 109125 118355 109191 118358
rect 113766 118356 113772 118420
rect 113836 118418 113842 118420
rect 253974 118418 253980 118420
rect 113836 118358 253980 118418
rect 113836 118356 113842 118358
rect 253974 118356 253980 118358
rect 254044 118418 254050 118420
rect 254853 118418 254919 118421
rect 254044 118416 254919 118418
rect 254044 118360 254858 118416
rect 254914 118360 254919 118416
rect 254044 118358 254919 118360
rect 254044 118356 254050 118358
rect 254853 118355 254919 118358
rect 5809 118282 5875 118285
rect 5809 118280 64890 118282
rect 5809 118224 5814 118280
rect 5870 118224 64890 118280
rect 5809 118222 64890 118224
rect 5809 118219 5875 118222
rect 55806 118084 55812 118148
rect 55876 118146 55882 118148
rect 56225 118146 56291 118149
rect 55876 118144 56291 118146
rect 55876 118088 56230 118144
rect 56286 118088 56291 118144
rect 55876 118086 56291 118088
rect 64830 118146 64890 118222
rect 79542 118220 79548 118284
rect 79612 118282 79618 118284
rect 168741 118282 168807 118285
rect 79612 118280 168807 118282
rect 79612 118224 168746 118280
rect 168802 118224 168807 118280
rect 79612 118222 168807 118224
rect 79612 118220 79618 118222
rect 168741 118219 168807 118222
rect 188981 118282 189047 118285
rect 205030 118282 205036 118284
rect 188981 118280 205036 118282
rect 188981 118224 188986 118280
rect 189042 118224 205036 118280
rect 188981 118222 205036 118224
rect 188981 118219 189047 118222
rect 205030 118220 205036 118222
rect 205100 118220 205106 118284
rect 223614 118220 223620 118284
rect 223684 118282 223690 118284
rect 241697 118282 241763 118285
rect 223684 118280 241763 118282
rect 223684 118224 241702 118280
rect 241758 118224 241763 118280
rect 223684 118222 241763 118224
rect 223684 118220 223690 118222
rect 241697 118219 241763 118222
rect 246246 118220 246252 118284
rect 246316 118282 246322 118284
rect 246316 118222 258090 118282
rect 246316 118220 246322 118222
rect 76373 118146 76439 118149
rect 84326 118146 84332 118148
rect 64830 118144 84332 118146
rect 64830 118088 76378 118144
rect 76434 118088 84332 118144
rect 64830 118086 84332 118088
rect 55876 118084 55882 118086
rect 56225 118083 56291 118086
rect 76373 118083 76439 118086
rect 84326 118084 84332 118086
rect 84396 118084 84402 118148
rect 103278 118084 103284 118148
rect 103348 118146 103354 118148
rect 141918 118146 141924 118148
rect 103348 118086 141924 118146
rect 103348 118084 103354 118086
rect 141918 118084 141924 118086
rect 141988 118146 141994 118148
rect 142337 118146 142403 118149
rect 141988 118144 142403 118146
rect 141988 118088 142342 118144
rect 142398 118088 142403 118144
rect 141988 118086 142403 118088
rect 141988 118084 141994 118086
rect 142337 118083 142403 118086
rect 208894 118084 208900 118148
rect 208964 118146 208970 118148
rect 209129 118146 209195 118149
rect 208964 118144 209195 118146
rect 208964 118088 209134 118144
rect 209190 118088 209195 118144
rect 208964 118086 209195 118088
rect 258030 118146 258090 118222
rect 268469 118146 268535 118149
rect 269062 118146 269068 118148
rect 258030 118144 269068 118146
rect 258030 118088 268474 118144
rect 268530 118088 269068 118144
rect 258030 118086 269068 118088
rect 208964 118084 208970 118086
rect 209129 118083 209195 118086
rect 268469 118083 268535 118086
rect 269062 118084 269068 118086
rect 269132 118084 269138 118148
rect 3693 118010 3759 118013
rect 223614 118010 223620 118012
rect 3693 118008 223620 118010
rect 3693 117952 3698 118008
rect 3754 117952 223620 118008
rect 3693 117950 223620 117952
rect 3693 117947 3759 117950
rect 223614 117948 223620 117950
rect 223684 117948 223690 118012
rect 248873 118010 248939 118013
rect 249006 118010 249012 118012
rect 248873 118008 249012 118010
rect 248873 117952 248878 118008
rect 248934 117952 249012 118008
rect 248873 117950 249012 117952
rect 248873 117947 248939 117950
rect 249006 117948 249012 117950
rect 249076 117948 249082 118012
rect 28758 117812 28764 117876
rect 28828 117874 28834 117876
rect 29729 117874 29795 117877
rect 28828 117872 35910 117874
rect 28828 117816 29734 117872
rect 29790 117816 35910 117872
rect 28828 117814 35910 117816
rect 28828 117812 28834 117814
rect 29729 117811 29795 117814
rect 35850 117738 35910 117814
rect 121310 117812 121316 117876
rect 121380 117874 121386 117876
rect 122189 117874 122255 117877
rect 121380 117872 122255 117874
rect 121380 117816 122194 117872
rect 122250 117816 122255 117872
rect 121380 117814 122255 117816
rect 121380 117812 121386 117814
rect 122189 117811 122255 117814
rect 283414 117738 283420 117740
rect 35850 117678 283420 117738
rect 283414 117676 283420 117678
rect 283484 117676 283490 117740
rect 293902 117676 293908 117740
rect 293972 117738 293978 117740
rect 295149 117738 295215 117741
rect 293972 117736 295215 117738
rect 293972 117680 295154 117736
rect 295210 117680 295215 117736
rect 293972 117678 295215 117680
rect 293972 117676 293978 117678
rect 295149 117675 295215 117678
rect 36486 117404 36492 117468
rect 36556 117466 36562 117468
rect 36629 117466 36695 117469
rect 36556 117464 36695 117466
rect 36556 117408 36634 117464
rect 36690 117408 36695 117464
rect 36556 117406 36695 117408
rect 36556 117404 36562 117406
rect 36629 117403 36695 117406
rect 49550 117404 49556 117468
rect 49620 117466 49626 117468
rect 49877 117466 49943 117469
rect 49620 117464 49943 117466
rect 49620 117408 49882 117464
rect 49938 117408 49943 117464
rect 49620 117406 49943 117408
rect 49620 117404 49626 117406
rect 49877 117403 49943 117406
rect 62614 117404 62620 117468
rect 62684 117466 62690 117468
rect 62757 117466 62823 117469
rect 62684 117464 62823 117466
rect 62684 117408 62762 117464
rect 62818 117408 62823 117464
rect 62684 117406 62823 117408
rect 62684 117404 62690 117406
rect 62757 117403 62823 117406
rect 82854 117404 82860 117468
rect 82924 117466 82930 117468
rect 82997 117466 83063 117469
rect 82924 117464 83063 117466
rect 82924 117408 83002 117464
rect 83058 117408 83063 117464
rect 82924 117406 83063 117408
rect 82924 117404 82930 117406
rect 82997 117403 83063 117406
rect 135846 117404 135852 117468
rect 135916 117466 135922 117468
rect 135989 117466 136055 117469
rect 135916 117464 136055 117466
rect 135916 117408 135994 117464
rect 136050 117408 136055 117464
rect 135916 117406 136055 117408
rect 135916 117404 135922 117406
rect 135989 117403 136055 117406
rect 149513 117466 149579 117469
rect 149830 117466 149836 117468
rect 149513 117464 149836 117466
rect 149513 117408 149518 117464
rect 149574 117408 149836 117464
rect 149513 117406 149836 117408
rect 149513 117403 149579 117406
rect 149830 117404 149836 117406
rect 149900 117404 149906 117468
rect 155350 117404 155356 117468
rect 155420 117466 155426 117468
rect 155585 117466 155651 117469
rect 155420 117464 155651 117466
rect 155420 117408 155590 117464
rect 155646 117408 155651 117464
rect 155420 117406 155651 117408
rect 155420 117404 155426 117406
rect 155585 117403 155651 117406
rect 161974 117404 161980 117468
rect 162044 117466 162050 117468
rect 162209 117466 162275 117469
rect 175917 117468 175983 117469
rect 175917 117466 175964 117468
rect 162044 117464 162275 117466
rect 162044 117408 162214 117464
rect 162270 117408 162275 117464
rect 162044 117406 162275 117408
rect 175872 117464 175964 117466
rect 175872 117408 175922 117464
rect 175872 117406 175964 117408
rect 162044 117404 162050 117406
rect 162209 117403 162275 117406
rect 175917 117404 175964 117406
rect 176028 117404 176034 117468
rect 182633 117466 182699 117469
rect 185158 117466 185164 117468
rect 182633 117464 185164 117466
rect 182633 117408 182638 117464
rect 182694 117408 185164 117464
rect 182633 117406 185164 117408
rect 175917 117403 175983 117404
rect 182633 117403 182699 117406
rect 185158 117404 185164 117406
rect 185228 117404 185234 117468
rect 188838 117404 188844 117468
rect 188908 117466 188914 117468
rect 188981 117466 189047 117469
rect 188908 117464 189047 117466
rect 188908 117408 188986 117464
rect 189042 117408 189047 117464
rect 188908 117406 189047 117408
rect 188908 117404 188914 117406
rect 188981 117403 189047 117406
rect 195094 117404 195100 117468
rect 195164 117466 195170 117468
rect 195329 117466 195395 117469
rect 195164 117464 195395 117466
rect 195164 117408 195334 117464
rect 195390 117408 195395 117464
rect 195164 117406 195395 117408
rect 195164 117404 195170 117406
rect 195329 117403 195395 117406
rect 202086 117404 202092 117468
rect 202156 117466 202162 117468
rect 202229 117466 202295 117469
rect 202156 117464 202295 117466
rect 202156 117408 202234 117464
rect 202290 117408 202295 117464
rect 202156 117406 202295 117408
rect 202156 117404 202162 117406
rect 202229 117403 202295 117406
rect 228214 117404 228220 117468
rect 228284 117466 228290 117468
rect 228817 117466 228883 117469
rect 228284 117464 228883 117466
rect 228284 117408 228822 117464
rect 228878 117408 228883 117464
rect 228284 117406 228883 117408
rect 228284 117404 228290 117406
rect 228817 117403 228883 117406
rect 235625 117466 235691 117469
rect 241697 117468 241763 117469
rect 235758 117466 235764 117468
rect 235625 117464 235764 117466
rect 235625 117408 235630 117464
rect 235686 117408 235764 117464
rect 235625 117406 235764 117408
rect 235625 117403 235691 117406
rect 235758 117404 235764 117406
rect 235828 117404 235834 117468
rect 241646 117404 241652 117468
rect 241716 117466 241763 117468
rect 281993 117466 282059 117469
rect 282126 117466 282132 117468
rect 241716 117464 241808 117466
rect 241758 117408 241808 117464
rect 241716 117406 241808 117408
rect 281993 117464 282132 117466
rect 281993 117408 281998 117464
rect 282054 117408 282132 117464
rect 281993 117406 282132 117408
rect 241716 117404 241763 117406
rect 241697 117403 241763 117404
rect 281993 117403 282059 117406
rect 282126 117404 282132 117406
rect 282196 117404 282202 117468
rect 3141 117330 3207 117333
rect 287094 117330 287100 117332
rect 3141 117328 287100 117330
rect 3141 117272 3146 117328
rect 3202 117272 287100 117328
rect 3141 117270 287100 117272
rect 3141 117267 3207 117270
rect 287094 117268 287100 117270
rect 287164 117330 287170 117332
rect 287973 117330 288039 117333
rect 287164 117328 288039 117330
rect 287164 117272 287978 117328
rect 288034 117272 288039 117328
rect 287164 117270 288039 117272
rect 287164 117268 287170 117270
rect 287973 117267 288039 117270
rect -960 116092 480 116332
rect 499520 116092 500960 116332
rect 209865 115834 209931 115837
rect 209998 115834 210004 115836
rect 209865 115832 210004 115834
rect 209865 115776 209870 115832
rect 209926 115776 210004 115832
rect 209865 115774 210004 115776
rect 209865 115771 209931 115774
rect 209998 115772 210004 115774
rect 210068 115772 210074 115836
rect 69381 114474 69447 114477
rect 70894 114474 70900 114476
rect 69381 114472 70900 114474
rect 69381 114416 69386 114472
rect 69442 114416 70900 114472
rect 69381 114414 70900 114416
rect 69381 114411 69447 114414
rect 70894 114412 70900 114414
rect 70964 114412 70970 114476
rect 7281 113930 7347 113933
rect 32489 113930 32555 113933
rect 303286 113930 303292 113932
rect 7281 113928 303292 113930
rect 7281 113872 7286 113928
rect 7342 113872 32494 113928
rect 32550 113872 303292 113928
rect 7281 113870 303292 113872
rect 7281 113867 7347 113870
rect 32489 113867 32555 113870
rect 303286 113868 303292 113870
rect 303356 113868 303362 113932
rect 186814 113052 186820 113116
rect 186884 113114 186890 113116
rect 187417 113114 187483 113117
rect 186884 113112 187483 113114
rect 186884 113056 187422 113112
rect 187478 113056 187483 113112
rect 186884 113054 187483 113056
rect 186884 113052 186890 113054
rect 187417 113051 187483 113054
rect 193070 113052 193076 113116
rect 193140 113114 193146 113116
rect 194041 113114 194107 113117
rect 193140 113112 194107 113114
rect 193140 113056 194046 113112
rect 194102 113056 194107 113112
rect 193140 113054 194107 113056
rect 193140 113052 193146 113054
rect 194041 113051 194107 113054
rect 219382 113052 219388 113116
rect 219452 113114 219458 113116
rect 220537 113114 220603 113117
rect 219452 113112 220603 113114
rect 219452 113056 220542 113112
rect 220598 113056 220603 113112
rect 219452 113054 220603 113056
rect 219452 113052 219458 113054
rect 220537 113051 220603 113054
rect 226926 113052 226932 113116
rect 226996 113114 227002 113116
rect 227161 113114 227227 113117
rect 226996 113112 227227 113114
rect 226996 113056 227166 113112
rect 227222 113056 227227 113112
rect 226996 113054 227227 113056
rect 226996 113052 227002 113054
rect 227161 113051 227227 113054
rect 273110 113052 273116 113116
rect 273180 113114 273186 113116
rect 273253 113114 273319 113117
rect 273180 113112 273319 113114
rect 273180 113056 273258 113112
rect 273314 113056 273319 113112
rect 273180 113054 273319 113056
rect 273180 113052 273186 113054
rect 273253 113051 273319 113054
rect 160921 112842 160987 112845
rect 162894 112842 162900 112844
rect 160921 112840 162900 112842
rect 160921 112784 160926 112840
rect 160982 112784 162900 112840
rect 160921 112782 162900 112784
rect 160921 112779 160987 112782
rect 162894 112780 162900 112782
rect 162964 112780 162970 112844
rect 167545 112842 167611 112845
rect 172462 112842 172468 112844
rect 167545 112840 172468 112842
rect 167545 112784 167550 112840
rect 167606 112784 172468 112840
rect 167545 112782 172468 112784
rect 167545 112779 167611 112782
rect 172462 112780 172468 112782
rect 172532 112780 172538 112844
rect 146886 112644 146892 112708
rect 146956 112706 146962 112708
rect 200665 112706 200731 112709
rect 146956 112704 200731 112706
rect 146956 112648 200670 112704
rect 200726 112648 200731 112704
rect 146956 112646 200731 112648
rect 146956 112644 146962 112646
rect 200665 112643 200731 112646
rect 213913 112706 213979 112709
rect 225086 112706 225092 112708
rect 213913 112704 225092 112706
rect 213913 112648 213918 112704
rect 213974 112648 225092 112704
rect 213913 112646 225092 112648
rect 213913 112643 213979 112646
rect 225086 112644 225092 112646
rect 225156 112644 225162 112708
rect 96654 112508 96660 112572
rect 96724 112570 96730 112572
rect 107929 112570 107995 112573
rect 96724 112568 107995 112570
rect 96724 112512 107934 112568
rect 107990 112512 107995 112568
rect 96724 112510 107995 112512
rect 96724 112508 96730 112510
rect 107929 112507 107995 112510
rect 141049 112570 141115 112573
rect 201534 112570 201540 112572
rect 141049 112568 201540 112570
rect 141049 112512 141054 112568
rect 141110 112512 201540 112568
rect 141049 112510 201540 112512
rect 141049 112507 141115 112510
rect 201534 112508 201540 112510
rect 201604 112508 201610 112572
rect 205950 112508 205956 112572
rect 206020 112570 206026 112572
rect 286777 112570 286843 112573
rect 206020 112568 286843 112570
rect 206020 112512 286782 112568
rect 286838 112512 286843 112568
rect 206020 112510 286843 112512
rect 206020 112508 206026 112510
rect 286777 112507 286843 112510
rect 149646 112372 149652 112436
rect 149716 112434 149722 112436
rect 247033 112434 247099 112437
rect 149716 112432 247099 112434
rect 149716 112376 247038 112432
rect 247094 112376 247099 112432
rect 149716 112374 247099 112376
rect 149716 112372 149722 112374
rect 247033 112371 247099 112374
rect 180793 112298 180859 112301
rect 184974 112298 184980 112300
rect 180793 112296 184980 112298
rect 180793 112240 180798 112296
rect 180854 112240 184980 112296
rect 180793 112238 184980 112240
rect 180793 112235 180859 112238
rect 184974 112236 184980 112238
rect 185044 112236 185050 112300
rect 52310 112100 52316 112164
rect 52380 112162 52386 112164
rect 52380 112102 55230 112162
rect 52380 112100 52386 112102
rect 9857 112026 9923 112029
rect 34462 112026 34468 112028
rect 9857 112024 34468 112026
rect -960 111740 480 111980
rect 9857 111968 9862 112024
rect 9918 111968 34468 112024
rect 9857 111966 34468 111968
rect 9857 111963 9923 111966
rect 34462 111964 34468 111966
rect 34532 112026 34538 112028
rect 35065 112026 35131 112029
rect 34532 112024 35131 112026
rect 34532 111968 35070 112024
rect 35126 111968 35131 112024
rect 34532 111966 35131 111968
rect 34532 111964 34538 111966
rect 35065 111963 35131 111966
rect 41689 112026 41755 112029
rect 42006 112026 42012 112028
rect 41689 112024 42012 112026
rect 41689 111968 41694 112024
rect 41750 111968 42012 112024
rect 41689 111966 42012 111968
rect 41689 111963 41755 111966
rect 42006 111964 42012 111966
rect 42076 111964 42082 112028
rect 54334 111964 54340 112028
rect 54404 112026 54410 112028
rect 54937 112026 55003 112029
rect 54404 112024 55003 112026
rect 54404 111968 54942 112024
rect 54998 111968 55003 112024
rect 54404 111966 55003 111968
rect 55170 112026 55230 112102
rect 59118 112100 59124 112164
rect 59188 112162 59194 112164
rect 61561 112162 61627 112165
rect 68185 112164 68251 112165
rect 115105 112164 115171 112165
rect 134425 112164 134491 112165
rect 59188 112160 61627 112162
rect 59188 112104 61566 112160
rect 61622 112104 61627 112160
rect 59188 112102 61627 112104
rect 59188 112100 59194 112102
rect 61561 112099 61627 112102
rect 68134 112100 68140 112164
rect 68204 112162 68251 112164
rect 115054 112162 115060 112164
rect 68204 112160 68296 112162
rect 68246 112104 68296 112160
rect 68204 112102 68296 112104
rect 115014 112102 115060 112162
rect 115124 112160 115171 112164
rect 115166 112104 115171 112160
rect 68204 112100 68251 112102
rect 115054 112100 115060 112102
rect 115124 112100 115171 112104
rect 134374 112100 134380 112164
rect 134444 112162 134491 112164
rect 134444 112160 134536 112162
rect 134486 112104 134536 112160
rect 134444 112102 134536 112104
rect 134444 112100 134491 112102
rect 145414 112100 145420 112164
rect 145484 112162 145490 112164
rect 147673 112162 147739 112165
rect 145484 112160 147739 112162
rect 145484 112104 147678 112160
rect 147734 112104 147739 112160
rect 145484 112102 147739 112104
rect 145484 112100 145490 112102
rect 68185 112099 68251 112100
rect 115105 112099 115171 112100
rect 134425 112099 134491 112100
rect 147673 112099 147739 112102
rect 153694 112100 153700 112164
rect 153764 112162 153770 112164
rect 154297 112162 154363 112165
rect 153764 112160 154363 112162
rect 153764 112104 154302 112160
rect 154358 112104 154363 112160
rect 153764 112102 154363 112104
rect 153764 112100 153770 112102
rect 154297 112099 154363 112102
rect 74809 112026 74875 112029
rect 83958 112026 83964 112028
rect 55170 112024 83964 112026
rect 55170 111968 74814 112024
rect 74870 111968 83964 112024
rect 55170 111966 83964 111968
rect 54404 111964 54410 111966
rect 54937 111963 55003 111966
rect 74809 111963 74875 111966
rect 83958 111964 83964 111966
rect 84028 111964 84034 112028
rect 87454 111964 87460 112028
rect 87524 112026 87530 112028
rect 88057 112026 88123 112029
rect 87524 112024 88123 112026
rect 87524 111968 88062 112024
rect 88118 111968 88123 112024
rect 87524 111966 88123 111968
rect 87524 111964 87530 111966
rect 88057 111963 88123 111966
rect 94446 111964 94452 112028
rect 94516 112026 94522 112028
rect 94681 112026 94747 112029
rect 101305 112028 101371 112029
rect 94516 112024 94747 112026
rect 94516 111968 94686 112024
rect 94742 111968 94747 112024
rect 94516 111966 94747 111968
rect 94516 111964 94522 111966
rect 94681 111963 94747 111966
rect 101254 111964 101260 112028
rect 101324 112026 101371 112028
rect 101324 112024 101416 112026
rect 101366 111968 101416 112024
rect 101324 111966 101416 111968
rect 101324 111964 101371 111966
rect 108430 111964 108436 112028
rect 108500 112026 108506 112028
rect 233785 112026 233851 112029
rect 108500 112024 234630 112026
rect 108500 111968 233790 112024
rect 233846 111968 234630 112024
rect 108500 111966 234630 111968
rect 108500 111964 108506 111966
rect 101305 111963 101371 111964
rect 233785 111963 233851 111966
rect 4061 111890 4127 111893
rect 173934 111890 173940 111892
rect 4061 111888 173940 111890
rect 4061 111832 4066 111888
rect 4122 111832 173940 111888
rect 4061 111830 173940 111832
rect 4061 111827 4127 111830
rect 173934 111828 173940 111830
rect 174004 111890 174010 111892
rect 174169 111890 174235 111893
rect 174004 111888 174235 111890
rect 174004 111832 174174 111888
rect 174230 111832 174235 111888
rect 174004 111830 174235 111832
rect 174004 111828 174010 111830
rect 174169 111827 174235 111830
rect 204110 111828 204116 111892
rect 204180 111890 204186 111892
rect 207289 111890 207355 111893
rect 204180 111888 207355 111890
rect 204180 111832 207294 111888
rect 207350 111832 207355 111888
rect 204180 111830 207355 111832
rect 234570 111890 234630 111966
rect 235942 111890 235948 111892
rect 234570 111830 235948 111890
rect 204180 111828 204186 111830
rect 207289 111827 207355 111830
rect 235942 111828 235948 111830
rect 236012 111828 236018 111892
rect 240174 111828 240180 111892
rect 240244 111890 240250 111892
rect 240409 111890 240475 111893
rect 240244 111888 240475 111890
rect 240244 111832 240414 111888
rect 240470 111832 240475 111888
rect 240244 111830 240475 111832
rect 240244 111828 240250 111830
rect 240409 111827 240475 111830
rect 253054 111828 253060 111892
rect 253124 111890 253130 111892
rect 253657 111890 253723 111893
rect 253124 111888 253723 111890
rect 253124 111832 253662 111888
rect 253718 111832 253723 111888
rect 253124 111830 253723 111832
rect 253124 111828 253130 111830
rect 253657 111827 253723 111830
rect 280153 111890 280219 111893
rect 280654 111890 280660 111892
rect 280153 111888 280660 111890
rect 280153 111832 280158 111888
rect 280214 111832 280660 111888
rect 280153 111830 280660 111832
rect 280153 111827 280219 111830
rect 280654 111828 280660 111830
rect 280724 111828 280730 111892
rect 293166 111828 293172 111892
rect 293236 111890 293242 111892
rect 293401 111890 293467 111893
rect 293236 111888 293467 111890
rect 293236 111832 293406 111888
rect 293462 111832 293467 111888
rect 293236 111830 293467 111832
rect 293236 111828 293242 111830
rect 293401 111827 293467 111830
rect 159214 111692 159220 111756
rect 159284 111754 159290 111756
rect 180609 111754 180675 111757
rect 159284 111752 180675 111754
rect 159284 111696 180614 111752
rect 180670 111696 180675 111752
rect 159284 111694 180675 111696
rect 159284 111692 159290 111694
rect 180609 111691 180675 111694
rect 132769 111620 132835 111621
rect 132718 111618 132724 111620
rect 132678 111558 132724 111618
rect 132788 111616 132835 111620
rect 132830 111560 132835 111616
rect 132718 111556 132724 111558
rect 132788 111556 132835 111560
rect 138606 111556 138612 111620
rect 138676 111618 138682 111620
rect 181253 111618 181319 111621
rect 138676 111616 181319 111618
rect 138676 111560 181258 111616
rect 181314 111560 181319 111616
rect 138676 111558 181319 111560
rect 138676 111556 138682 111558
rect 132769 111555 132835 111556
rect 181253 111555 181319 111558
rect 130326 111420 130332 111484
rect 130396 111482 130402 111484
rect 179505 111482 179571 111485
rect 130396 111480 179571 111482
rect 130396 111424 179510 111480
rect 179566 111424 179571 111480
rect 130396 111422 179571 111424
rect 130396 111420 130402 111422
rect 179505 111419 179571 111422
rect 213126 111420 213132 111484
rect 213196 111482 213202 111484
rect 213637 111482 213703 111485
rect 213196 111480 213703 111482
rect 213196 111424 213642 111480
rect 213698 111424 213703 111480
rect 499520 111468 500960 111708
rect 213196 111422 213703 111424
rect 213196 111420 213202 111422
rect 213637 111419 213703 111422
rect 128854 111284 128860 111348
rect 128924 111346 128930 111348
rect 179321 111346 179387 111349
rect 128924 111344 179387 111346
rect 128924 111288 179326 111344
rect 179382 111288 179387 111344
rect 128924 111286 179387 111288
rect 128924 111284 128930 111286
rect 179321 111283 179387 111286
rect 182633 111346 182699 111349
rect 183461 111346 183527 111349
rect 182633 111344 183527 111346
rect 182633 111288 182638 111344
rect 182694 111288 183466 111344
rect 183522 111288 183527 111344
rect 182633 111286 183527 111288
rect 182633 111283 182699 111286
rect 183461 111283 183527 111286
rect 188286 111284 188292 111348
rect 188356 111346 188362 111348
rect 214465 111346 214531 111349
rect 188356 111344 214531 111346
rect 188356 111288 214470 111344
rect 214526 111288 214531 111344
rect 188356 111286 214531 111288
rect 188356 111284 188362 111286
rect 214465 111283 214531 111286
rect 111006 111148 111012 111212
rect 111076 111210 111082 111212
rect 170213 111210 170279 111213
rect 111076 111208 170279 111210
rect 111076 111152 170218 111208
rect 170274 111152 170279 111208
rect 111076 111150 170279 111152
rect 111076 111148 111082 111150
rect 170213 111147 170279 111150
rect 181805 111210 181871 111213
rect 183185 111210 183251 111213
rect 181805 111208 183251 111210
rect 181805 111152 181810 111208
rect 181866 111152 183190 111208
rect 183246 111152 183251 111208
rect 181805 111150 183251 111152
rect 181805 111147 181871 111150
rect 183185 111147 183251 111150
rect 191046 111148 191052 111212
rect 191116 111210 191122 111212
rect 222377 111210 222443 111213
rect 191116 111208 222443 111210
rect 191116 111152 222382 111208
rect 222438 111152 222443 111208
rect 191116 111150 222443 111152
rect 191116 111148 191122 111150
rect 222377 111147 222443 111150
rect 231853 111210 231919 111213
rect 232446 111210 232452 111212
rect 231853 111208 232452 111210
rect 231853 111152 231858 111208
rect 231914 111152 232452 111208
rect 231853 111150 232452 111152
rect 231853 111147 231919 111150
rect 232446 111148 232452 111150
rect 232516 111148 232522 111212
rect 124806 111012 124812 111076
rect 124876 111074 124882 111076
rect 194409 111074 194475 111077
rect 124876 111072 194475 111074
rect 124876 111016 194414 111072
rect 194470 111016 194475 111072
rect 124876 111014 194475 111016
rect 124876 111012 124882 111014
rect 194409 111011 194475 111014
rect 214649 111074 214715 111077
rect 274030 111074 274036 111076
rect 214649 111072 274036 111074
rect 214649 111016 214654 111072
rect 214710 111016 274036 111072
rect 214649 111014 274036 111016
rect 214649 111011 214715 111014
rect 274030 111012 274036 111014
rect 274100 111012 274106 111076
rect 135713 110938 135779 110941
rect 214557 110938 214623 110941
rect 135713 110936 214623 110938
rect 135713 110880 135718 110936
rect 135774 110880 214562 110936
rect 214618 110880 214623 110936
rect 135713 110878 214623 110880
rect 135713 110875 135779 110878
rect 214557 110875 214623 110878
rect 214741 110938 214807 110941
rect 220854 110938 220860 110940
rect 214741 110936 220860 110938
rect 214741 110880 214746 110936
rect 214802 110880 220860 110936
rect 214741 110878 220860 110880
rect 214741 110875 214807 110878
rect 220854 110876 220860 110878
rect 220924 110876 220930 110940
rect 51574 110740 51580 110804
rect 51644 110802 51650 110804
rect 168373 110802 168439 110805
rect 51644 110800 168439 110802
rect 51644 110744 168378 110800
rect 168434 110744 168439 110800
rect 51644 110742 168439 110744
rect 51644 110740 51650 110742
rect 168373 110739 168439 110742
rect 175774 110740 175780 110804
rect 175844 110802 175850 110804
rect 273805 110802 273871 110805
rect 175844 110800 273871 110802
rect 175844 110744 273810 110800
rect 273866 110744 273871 110800
rect 175844 110742 273871 110744
rect 175844 110740 175850 110742
rect 273805 110739 273871 110742
rect 90766 110604 90772 110668
rect 90836 110666 90842 110668
rect 96889 110666 96955 110669
rect 90836 110664 96955 110666
rect 90836 110608 96894 110664
rect 96950 110608 96955 110664
rect 90836 110606 96955 110608
rect 90836 110604 90842 110606
rect 96889 110603 96955 110606
rect 108246 110604 108252 110668
rect 108316 110666 108322 110668
rect 273161 110666 273227 110669
rect 108316 110664 273227 110666
rect 108316 110608 273166 110664
rect 273222 110608 273227 110664
rect 108316 110606 273227 110608
rect 108316 110604 108322 110606
rect 273161 110603 273227 110606
rect 137185 110530 137251 110533
rect 138790 110530 138796 110532
rect 137185 110528 138796 110530
rect 137185 110472 137190 110528
rect 137246 110472 138796 110528
rect 137185 110470 138796 110472
rect 137185 110467 137251 110470
rect 138790 110468 138796 110470
rect 138860 110468 138866 110532
rect 155166 110468 155172 110532
rect 155236 110530 155242 110532
rect 168097 110530 168163 110533
rect 182633 110532 182699 110533
rect 182582 110530 182588 110532
rect 155236 110528 168163 110530
rect 155236 110472 168102 110528
rect 168158 110472 168163 110528
rect 155236 110470 168163 110472
rect 182542 110470 182588 110530
rect 182652 110528 182699 110532
rect 182694 110472 182699 110528
rect 155236 110468 155242 110470
rect 168097 110467 168163 110470
rect 182582 110468 182588 110470
rect 182652 110468 182699 110472
rect 182633 110467 182699 110468
rect 190453 110532 190519 110533
rect 190453 110528 190500 110532
rect 190564 110530 190570 110532
rect 190453 110472 190458 110528
rect 190453 110468 190500 110472
rect 190564 110470 190610 110530
rect 190564 110468 190570 110470
rect 209078 110468 209084 110532
rect 209148 110530 209154 110532
rect 222193 110530 222259 110533
rect 273621 110532 273687 110533
rect 222326 110530 222332 110532
rect 209148 110528 222332 110530
rect 209148 110472 222198 110528
rect 222254 110472 222332 110528
rect 209148 110470 222332 110472
rect 209148 110468 209154 110470
rect 190453 110467 190519 110468
rect 222193 110467 222259 110470
rect 222326 110468 222332 110470
rect 222396 110468 222402 110532
rect 273621 110528 273668 110532
rect 273732 110530 273738 110532
rect 273621 110472 273626 110528
rect 273621 110468 273668 110472
rect 273732 110470 273778 110530
rect 273732 110468 273738 110470
rect 273621 110467 273687 110468
rect 88149 109444 88215 109445
rect 88149 109442 88196 109444
rect 88104 109440 88196 109442
rect 88104 109384 88154 109440
rect 88104 109382 88196 109384
rect 88149 109380 88196 109382
rect 88260 109380 88266 109444
rect 88149 109379 88215 109380
rect 9121 109170 9187 109173
rect 293902 109170 293908 109172
rect 9121 109168 293908 109170
rect 9121 109112 9126 109168
rect 9182 109112 293908 109168
rect 9121 109110 293908 109112
rect 9121 109107 9187 109110
rect 293902 109108 293908 109110
rect 293972 109108 293978 109172
rect 7925 108626 7991 108629
rect 7925 108624 10058 108626
rect 7925 108568 7930 108624
rect 7986 108568 10058 108624
rect 7925 108566 10058 108568
rect 7925 108563 7991 108566
rect 9998 107984 10058 108566
rect 81934 108292 81940 108356
rect 82004 108354 82010 108356
rect 182582 108354 182588 108356
rect 82004 108294 182588 108354
rect 82004 108292 82010 108294
rect 182582 108292 182588 108294
rect 182652 108292 182658 108356
rect -960 107388 480 107628
rect 499520 107116 500960 107356
rect 312629 105634 312695 105637
rect 309918 105632 312695 105634
rect 309918 105576 312634 105632
rect 312690 105576 312695 105632
rect 309918 105574 312695 105576
rect 309918 104992 309978 105574
rect 312629 105571 312695 105574
rect -960 102764 480 103004
rect 495525 102642 495591 102645
rect 499520 102642 500960 102732
rect 495525 102640 500960 102642
rect 495525 102584 495530 102640
rect 495586 102584 500960 102640
rect 495525 102582 500960 102584
rect 495525 102579 495591 102582
rect 499520 102492 500960 102582
rect 8017 98834 8083 98837
rect 8017 98832 10058 98834
rect 8017 98776 8022 98832
rect 8078 98776 10058 98832
rect 8017 98774 10058 98776
rect 8017 98771 8083 98774
rect -960 98412 480 98652
rect 9998 98192 10058 98774
rect 495525 98290 495591 98293
rect 499520 98290 500960 98380
rect 495525 98288 500960 98290
rect 495525 98232 495530 98288
rect 495586 98232 500960 98288
rect 495525 98230 500960 98232
rect 495525 98227 495591 98230
rect 499520 98140 500960 98230
rect 309918 95162 309978 95200
rect 312537 95162 312603 95165
rect 309918 95160 312603 95162
rect 309918 95104 312542 95160
rect 312598 95104 312603 95160
rect 309918 95102 312603 95104
rect 312537 95099 312603 95102
rect -960 93788 480 94028
rect 495525 93666 495591 93669
rect 499520 93666 500960 93756
rect 495525 93664 500960 93666
rect 495525 93608 495530 93664
rect 495586 93608 500960 93664
rect 495525 93606 500960 93608
rect 495525 93603 495591 93606
rect 499520 93516 500960 93606
rect -960 89436 480 89676
rect 495525 89314 495591 89317
rect 499520 89314 500960 89404
rect 495525 89312 500960 89314
rect 495525 89256 495530 89312
rect 495586 89256 500960 89312
rect 495525 89254 500960 89256
rect 495525 89251 495591 89254
rect 499520 89164 500960 89254
rect 8017 89042 8083 89045
rect 8017 89040 10058 89042
rect 8017 88984 8022 89040
rect 8078 88984 10058 89040
rect 8017 88982 10058 88984
rect 8017 88979 8083 88982
rect 9998 88400 10058 88982
rect 311985 85506 312051 85509
rect 309918 85504 312051 85506
rect 309918 85448 311990 85504
rect 312046 85448 312051 85504
rect 309918 85446 312051 85448
rect 309918 85408 309978 85446
rect 311985 85443 312051 85446
rect -960 84962 480 85052
rect 3785 84962 3851 84965
rect -960 84960 3851 84962
rect -960 84904 3790 84960
rect 3846 84904 3851 84960
rect -960 84902 3851 84904
rect -960 84812 480 84902
rect 3785 84899 3851 84902
rect 499520 84540 500960 84780
rect -960 80610 480 80700
rect 3509 80610 3575 80613
rect -960 80608 3575 80610
rect -960 80552 3514 80608
rect 3570 80552 3575 80608
rect -960 80550 3575 80552
rect -960 80460 480 80550
rect 3509 80547 3575 80550
rect 499520 80188 500960 80428
rect 8109 78570 8175 78573
rect 9998 78570 10058 78608
rect 8109 78568 10058 78570
rect 8109 78512 8114 78568
rect 8170 78512 10058 78568
rect 8109 78510 10058 78512
rect 8109 78507 8175 78510
rect -960 75986 480 76076
rect 2773 75986 2839 75989
rect -960 75984 2839 75986
rect -960 75928 2778 75984
rect 2834 75928 2839 75984
rect -960 75926 2839 75928
rect -960 75836 480 75926
rect 2773 75923 2839 75926
rect 312445 75850 312511 75853
rect 309918 75848 312511 75850
rect 309918 75792 312450 75848
rect 312506 75792 312511 75848
rect 309918 75790 312511 75792
rect 309918 75616 309978 75790
rect 312445 75787 312511 75790
rect 499520 75564 500960 75804
rect -960 71484 480 71724
rect 499520 71212 500960 71452
rect 7465 68914 7531 68917
rect 7465 68912 10058 68914
rect 7465 68856 7470 68912
rect 7526 68856 10058 68912
rect 7465 68854 10058 68856
rect 7465 68851 7531 68854
rect 9998 68816 10058 68854
rect -960 67010 480 67100
rect 3141 67010 3207 67013
rect -960 67008 3207 67010
rect -960 66952 3146 67008
rect 3202 66952 3207 67008
rect -960 66950 3207 66952
rect -960 66860 480 66950
rect 3141 66947 3207 66950
rect 499520 66860 500960 67100
rect 312353 66194 312419 66197
rect 309918 66192 312419 66194
rect 309918 66136 312358 66192
rect 312414 66136 312419 66192
rect 309918 66134 312419 66136
rect 309918 65824 309978 66134
rect 312353 66131 312419 66134
rect -960 62508 480 62748
rect 495525 62386 495591 62389
rect 499520 62386 500960 62476
rect 495525 62384 500960 62386
rect 495525 62328 495530 62384
rect 495586 62328 500960 62384
rect 495525 62326 500960 62328
rect 495525 62323 495591 62326
rect 499520 62236 500960 62326
rect 7373 59258 7439 59261
rect 8109 59258 8175 59261
rect 7373 59256 10058 59258
rect 7373 59200 7378 59256
rect 7434 59200 8114 59256
rect 8170 59200 10058 59256
rect 7373 59198 10058 59200
rect 7373 59195 7439 59198
rect 8109 59195 8175 59198
rect 9998 59024 10058 59198
rect -960 58034 480 58124
rect 2773 58034 2839 58037
rect -960 58032 2839 58034
rect -960 57976 2778 58032
rect 2834 57976 2839 58032
rect -960 57974 2839 57976
rect -960 57884 480 57974
rect 2773 57971 2839 57974
rect 495525 58034 495591 58037
rect 499520 58034 500960 58124
rect 495525 58032 500960 58034
rect 495525 57976 495530 58032
rect 495586 57976 500960 58032
rect 495525 57974 500960 57976
rect 495525 57971 495591 57974
rect 499520 57884 500960 57974
rect 309918 55994 309978 56032
rect 312077 55994 312143 55997
rect 312445 55994 312511 55997
rect 309918 55992 312511 55994
rect 309918 55936 312082 55992
rect 312138 55936 312450 55992
rect 312506 55936 312511 55992
rect 309918 55934 312511 55936
rect 312077 55931 312143 55934
rect 312445 55931 312511 55934
rect -960 53682 480 53772
rect 2773 53682 2839 53685
rect -960 53680 2839 53682
rect -960 53624 2778 53680
rect 2834 53624 2839 53680
rect -960 53622 2839 53624
rect -960 53532 480 53622
rect 2773 53619 2839 53622
rect 499520 53260 500960 53500
rect 7189 49602 7255 49605
rect 7189 49600 10058 49602
rect 7189 49544 7194 49600
rect 7250 49544 10058 49600
rect 7189 49542 10058 49544
rect 7189 49539 7255 49542
rect -960 49180 480 49420
rect 9998 49232 10058 49542
rect 499520 48908 500960 49148
rect 309918 45930 309978 46240
rect 310605 45930 310671 45933
rect 309918 45928 310671 45930
rect 309918 45872 310610 45928
rect 310666 45872 310671 45928
rect 309918 45870 310671 45872
rect 310605 45867 310671 45870
rect -960 44706 480 44796
rect 4061 44706 4127 44709
rect -960 44704 4127 44706
rect -960 44648 4066 44704
rect 4122 44648 4127 44704
rect -960 44646 4127 44648
rect -960 44556 480 44646
rect 4061 44643 4127 44646
rect 495525 44434 495591 44437
rect 499520 44434 500960 44524
rect 495525 44432 500960 44434
rect 495525 44376 495530 44432
rect 495586 44376 500960 44432
rect 495525 44374 500960 44376
rect 495525 44371 495591 44374
rect 499520 44284 500960 44374
rect -960 40354 480 40444
rect 3233 40354 3299 40357
rect -960 40352 3299 40354
rect -960 40296 3238 40352
rect 3294 40296 3299 40352
rect -960 40294 3299 40296
rect -960 40204 480 40294
rect 3233 40291 3299 40294
rect 496169 40082 496235 40085
rect 499520 40082 500960 40172
rect 496169 40080 500960 40082
rect 496169 40024 496174 40080
rect 496230 40024 500960 40080
rect 496169 40022 500960 40024
rect 496169 40019 496235 40022
rect 7557 39946 7623 39949
rect 7557 39944 10058 39946
rect 7557 39888 7562 39944
rect 7618 39888 10058 39944
rect 499520 39932 500960 40022
rect 7557 39886 10058 39888
rect 7557 39883 7623 39886
rect 9998 39440 10058 39886
rect 312721 36682 312787 36685
rect 309918 36680 312787 36682
rect 309918 36624 312726 36680
rect 312782 36624 312787 36680
rect 309918 36622 312787 36624
rect 309918 36448 309978 36622
rect 312721 36619 312787 36622
rect -960 35730 480 35820
rect 3417 35730 3483 35733
rect -960 35728 3483 35730
rect -960 35672 3422 35728
rect 3478 35672 3483 35728
rect -960 35670 3483 35672
rect -960 35580 480 35670
rect 3417 35667 3483 35670
rect 495525 35458 495591 35461
rect 499520 35458 500960 35548
rect 495525 35456 500960 35458
rect 495525 35400 495530 35456
rect 495586 35400 500960 35456
rect 495525 35398 500960 35400
rect 495525 35395 495591 35398
rect 499520 35308 500960 35398
rect -960 31228 480 31468
rect 499520 30956 500960 31196
rect 7649 30290 7715 30293
rect 7649 30288 10058 30290
rect 7649 30232 7654 30288
rect 7710 30232 10058 30288
rect 7649 30230 10058 30232
rect 7649 30227 7715 30230
rect 9998 29648 10058 30230
rect 312537 27298 312603 27301
rect 309918 27296 312603 27298
rect 309918 27240 312542 27296
rect 312598 27240 312603 27296
rect 309918 27238 312603 27240
rect -960 26604 480 26844
rect 309918 26656 309978 27238
rect 312537 27235 312603 27238
rect 499520 26332 500960 26572
rect -960 22252 480 22492
rect 495525 22130 495591 22133
rect 499520 22130 500960 22220
rect 495525 22128 500960 22130
rect 495525 22072 495530 22128
rect 495586 22072 500960 22128
rect 495525 22070 500960 22072
rect 495525 22067 495591 22070
rect 499520 21980 500960 22070
rect 8201 20498 8267 20501
rect 8201 20496 10058 20498
rect 8201 20440 8206 20496
rect 8262 20440 10058 20496
rect 8201 20438 10058 20440
rect 8201 20435 8267 20438
rect 9998 19856 10058 20438
rect 311893 17914 311959 17917
rect 312261 17914 312327 17917
rect 311893 17912 312327 17914
rect -960 17778 480 17868
rect 311893 17856 311898 17912
rect 311954 17856 312266 17912
rect 312322 17856 312327 17912
rect 311893 17854 312327 17856
rect 311893 17851 311959 17854
rect 312261 17851 312327 17854
rect 3417 17778 3483 17781
rect -960 17776 3483 17778
rect -960 17720 3422 17776
rect 3478 17720 3483 17776
rect -960 17718 3483 17720
rect -960 17628 480 17718
rect 3417 17715 3483 17718
rect 499520 17356 500960 17596
rect 311893 16962 311959 16965
rect 309918 16960 311959 16962
rect 309918 16904 311898 16960
rect 311954 16904 311959 16960
rect 309918 16902 311959 16904
rect 309918 16864 309978 16902
rect 311893 16899 311959 16902
rect -960 13276 480 13516
rect 495433 13154 495499 13157
rect 499520 13154 500960 13244
rect 495433 13152 500960 13154
rect 495433 13096 495438 13152
rect 495494 13096 500960 13152
rect 495433 13094 500960 13096
rect 495433 13091 495499 13094
rect 499520 13004 500960 13094
rect 28758 10644 28764 10708
rect 28828 10706 28834 10708
rect 29637 10706 29703 10709
rect 28828 10704 29703 10706
rect 28828 10648 29642 10704
rect 29698 10648 29703 10704
rect 28828 10646 29703 10648
rect 28828 10644 28834 10646
rect 29637 10643 29703 10646
rect 49550 10644 49556 10708
rect 49620 10706 49626 10708
rect 49877 10706 49943 10709
rect 49620 10704 49943 10706
rect 49620 10648 49882 10704
rect 49938 10648 49943 10704
rect 49620 10646 49943 10648
rect 49620 10644 49626 10646
rect 49877 10643 49943 10646
rect 55806 10644 55812 10708
rect 55876 10706 55882 10708
rect 56133 10706 56199 10709
rect 55876 10704 56199 10706
rect 55876 10648 56138 10704
rect 56194 10648 56199 10704
rect 55876 10646 56199 10648
rect 55876 10644 55882 10646
rect 56133 10643 56199 10646
rect 62614 10644 62620 10708
rect 62684 10706 62690 10708
rect 62757 10706 62823 10709
rect 62684 10704 62823 10706
rect 62684 10648 62762 10704
rect 62818 10648 62823 10704
rect 62684 10646 62823 10648
rect 62684 10644 62690 10646
rect 62757 10643 62823 10646
rect 121310 10644 121316 10708
rect 121380 10706 121386 10708
rect 122373 10706 122439 10709
rect 121380 10704 122439 10706
rect 121380 10648 122378 10704
rect 122434 10648 122439 10704
rect 121380 10646 122439 10648
rect 121380 10644 121386 10646
rect 122373 10643 122439 10646
rect 155350 10644 155356 10708
rect 155420 10706 155426 10708
rect 155493 10706 155559 10709
rect 155420 10704 155559 10706
rect 155420 10648 155498 10704
rect 155554 10648 155559 10704
rect 155420 10646 155559 10648
rect 155420 10644 155426 10646
rect 155493 10643 155559 10646
rect 161974 10644 161980 10708
rect 162044 10706 162050 10708
rect 162117 10706 162183 10709
rect 175917 10708 175983 10709
rect 175917 10706 175964 10708
rect 162044 10704 162183 10706
rect 162044 10648 162122 10704
rect 162178 10648 162183 10704
rect 162044 10646 162183 10648
rect 175872 10704 175964 10706
rect 175872 10648 175922 10704
rect 175872 10646 175964 10648
rect 162044 10644 162050 10646
rect 162117 10643 162183 10646
rect 175917 10644 175964 10646
rect 176028 10644 176034 10708
rect 182633 10706 182699 10709
rect 185158 10706 185164 10708
rect 182633 10704 185164 10706
rect 182633 10648 182638 10704
rect 182694 10648 185164 10704
rect 182633 10646 185164 10648
rect 175917 10643 175983 10644
rect 182633 10643 182699 10646
rect 185158 10644 185164 10646
rect 185228 10644 185234 10708
rect 188838 10644 188844 10708
rect 188908 10706 188914 10708
rect 188981 10706 189047 10709
rect 188908 10704 189047 10706
rect 188908 10648 188986 10704
rect 189042 10648 189047 10704
rect 188908 10646 189047 10648
rect 188908 10644 188914 10646
rect 188981 10643 189047 10646
rect 195094 10644 195100 10708
rect 195164 10706 195170 10708
rect 195237 10706 195303 10709
rect 195164 10704 195303 10706
rect 195164 10648 195242 10704
rect 195298 10648 195303 10704
rect 195164 10646 195303 10648
rect 195164 10644 195170 10646
rect 195237 10643 195303 10646
rect 202086 10644 202092 10708
rect 202156 10706 202162 10708
rect 202229 10706 202295 10709
rect 208853 10708 208919 10709
rect 208853 10706 208900 10708
rect 202156 10704 202295 10706
rect 202156 10648 202234 10704
rect 202290 10648 202295 10704
rect 202156 10646 202295 10648
rect 208808 10704 208900 10706
rect 208808 10648 208858 10704
rect 208808 10646 208900 10648
rect 202156 10644 202162 10646
rect 202229 10643 202295 10646
rect 208853 10644 208900 10646
rect 208964 10644 208970 10708
rect 228214 10644 228220 10708
rect 228284 10706 228290 10708
rect 228357 10706 228423 10709
rect 228284 10704 228423 10706
rect 228284 10648 228362 10704
rect 228418 10648 228423 10704
rect 228284 10646 228423 10648
rect 228284 10644 228290 10646
rect 208853 10643 208919 10644
rect 228357 10643 228423 10646
rect 235625 10706 235691 10709
rect 235758 10706 235764 10708
rect 235625 10704 235764 10706
rect 235625 10648 235630 10704
rect 235686 10648 235764 10704
rect 235625 10646 235764 10648
rect 235625 10643 235691 10646
rect 235758 10644 235764 10646
rect 235828 10644 235834 10708
rect 248873 10706 248939 10709
rect 249006 10706 249012 10708
rect 248873 10704 249012 10706
rect 248873 10648 248878 10704
rect 248934 10648 249012 10704
rect 248873 10646 249012 10648
rect 248873 10643 248939 10646
rect 249006 10644 249012 10646
rect 249076 10644 249082 10708
rect 253974 10644 253980 10708
rect 254044 10706 254050 10708
rect 254853 10706 254919 10709
rect 254044 10704 254919 10706
rect 254044 10648 254858 10704
rect 254914 10648 254919 10704
rect 254044 10646 254919 10648
rect 254044 10644 254050 10646
rect 254853 10643 254919 10646
rect 261334 10644 261340 10708
rect 261404 10706 261410 10708
rect 261477 10706 261543 10709
rect 261404 10704 261543 10706
rect 261404 10648 261482 10704
rect 261538 10648 261543 10704
rect 261404 10646 261543 10648
rect 261404 10644 261410 10646
rect 261477 10643 261543 10646
rect 268745 10706 268811 10709
rect 269062 10706 269068 10708
rect 268745 10704 269068 10706
rect 268745 10648 268750 10704
rect 268806 10648 269068 10704
rect 268745 10646 269068 10648
rect 268745 10643 268811 10646
rect 269062 10644 269068 10646
rect 269132 10644 269138 10708
rect 273662 10644 273668 10708
rect 273732 10706 273738 10708
rect 274725 10706 274791 10709
rect 273732 10704 274791 10706
rect 273732 10648 274730 10704
rect 274786 10648 274791 10704
rect 273732 10646 274791 10648
rect 273732 10644 273738 10646
rect 274725 10643 274791 10646
rect 281993 10706 282059 10709
rect 282126 10706 282132 10708
rect 281993 10704 282132 10706
rect 281993 10648 281998 10704
rect 282054 10648 282132 10704
rect 281993 10646 282132 10648
rect 281993 10643 282059 10646
rect 282126 10644 282132 10646
rect 282196 10644 282202 10708
rect 287094 10644 287100 10708
rect 287164 10706 287170 10708
rect 287973 10706 288039 10709
rect 287164 10704 288039 10706
rect 287164 10648 287978 10704
rect 288034 10648 288039 10704
rect 287164 10646 288039 10648
rect 287164 10644 287170 10646
rect 287973 10643 288039 10646
rect 293902 10644 293908 10708
rect 293972 10706 293978 10708
rect 294597 10706 294663 10709
rect 293972 10704 294663 10706
rect 293972 10648 294602 10704
rect 294658 10648 294663 10704
rect 293972 10646 294663 10648
rect 293972 10644 293978 10646
rect 294597 10643 294663 10646
rect 215886 10236 215892 10300
rect 215956 10298 215962 10300
rect 244549 10298 244615 10301
rect 215956 10296 244615 10298
rect 215956 10240 244554 10296
rect 244610 10240 244615 10296
rect 215956 10238 244615 10240
rect 215956 10236 215962 10238
rect 244549 10235 244615 10238
rect 149513 10162 149579 10165
rect 241697 10164 241763 10165
rect 149830 10162 149836 10164
rect 149513 10160 149836 10162
rect 149513 10104 149518 10160
rect 149574 10104 149836 10160
rect 149513 10102 149836 10104
rect 149513 10099 149579 10102
rect 149830 10100 149836 10102
rect 149900 10100 149906 10164
rect 241646 10162 241652 10164
rect 241606 10102 241652 10162
rect 241716 10160 241763 10164
rect 241758 10104 241763 10160
rect 241646 10100 241652 10102
rect 241716 10100 241763 10104
rect 241697 10099 241763 10100
rect 36537 9892 36603 9893
rect 82905 9892 82971 9893
rect 135897 9892 135963 9893
rect 36486 9890 36492 9892
rect 36446 9830 36492 9890
rect 36556 9888 36603 9892
rect 82854 9890 82860 9892
rect 36598 9832 36603 9888
rect 36486 9828 36492 9830
rect 36556 9828 36603 9832
rect 82814 9830 82860 9890
rect 82924 9888 82971 9892
rect 135846 9890 135852 9892
rect 82966 9832 82971 9888
rect 82854 9828 82860 9830
rect 82924 9828 82971 9832
rect 135806 9830 135852 9890
rect 135916 9888 135963 9892
rect 135958 9832 135963 9888
rect 135846 9828 135852 9830
rect 135916 9828 135963 9832
rect 142102 9828 142108 9892
rect 142172 9890 142178 9892
rect 142245 9890 142311 9893
rect 142172 9888 142311 9890
rect 142172 9832 142250 9888
rect 142306 9832 142311 9888
rect 142172 9830 142311 9832
rect 142172 9828 142178 9830
rect 36537 9827 36603 9828
rect 82905 9827 82971 9828
rect 135897 9827 135963 9828
rect 142245 9827 142311 9830
rect 168465 9754 168531 9757
rect 168925 9754 168991 9757
rect 168465 9752 168991 9754
rect 168465 9696 168470 9752
rect 168526 9696 168930 9752
rect 168986 9696 168991 9752
rect 168465 9694 168991 9696
rect 168465 9691 168531 9694
rect 168925 9691 168991 9694
rect 69606 9556 69612 9620
rect 69676 9618 69682 9620
rect 77293 9618 77359 9621
rect 77845 9620 77911 9621
rect 77845 9618 77892 9620
rect 69676 9616 77359 9618
rect 69676 9560 77298 9616
rect 77354 9560 77359 9616
rect 69676 9558 77359 9560
rect 77800 9616 77892 9618
rect 77800 9560 77850 9616
rect 77800 9558 77892 9560
rect 69676 9556 69682 9558
rect 77293 9555 77359 9558
rect 77845 9556 77892 9558
rect 77956 9556 77962 9620
rect 78581 9618 78647 9621
rect 88926 9618 88932 9620
rect 78581 9616 88932 9618
rect 78581 9560 78586 9616
rect 78642 9560 88932 9616
rect 78581 9558 88932 9560
rect 77845 9555 77911 9556
rect 78581 9555 78647 9558
rect 88926 9556 88932 9558
rect 88996 9556 89002 9620
rect 95141 9618 95207 9621
rect 105486 9618 105492 9620
rect 95141 9616 105492 9618
rect 95141 9560 95146 9616
rect 95202 9560 105492 9616
rect 95141 9558 105492 9560
rect 95141 9555 95207 9558
rect 105486 9556 105492 9558
rect 105556 9556 105562 9620
rect 116485 9618 116551 9621
rect 117814 9618 117820 9620
rect 116485 9616 117820 9618
rect 116485 9560 116490 9616
rect 116546 9560 117820 9616
rect 116485 9558 117820 9560
rect 116485 9555 116551 9558
rect 117814 9556 117820 9558
rect 117884 9556 117890 9620
rect 168741 9618 168807 9621
rect 169293 9618 169359 9621
rect 168741 9616 169359 9618
rect 168741 9560 168746 9616
rect 168802 9560 169298 9616
rect 169354 9560 169359 9616
rect 168741 9558 169359 9560
rect 168741 9555 168807 9558
rect 169293 9555 169359 9558
rect 184054 9556 184060 9620
rect 184124 9618 184130 9620
rect 185761 9618 185827 9621
rect 272057 9618 272123 9621
rect 273161 9618 273227 9621
rect 184124 9616 185827 9618
rect 184124 9560 185766 9616
rect 185822 9560 185827 9616
rect 184124 9558 185827 9560
rect 184124 9556 184130 9558
rect 185761 9555 185827 9558
rect 238710 9558 253950 9618
rect 9121 9482 9187 9485
rect 65149 9482 65215 9485
rect 66161 9482 66227 9485
rect 9121 9480 66227 9482
rect 9121 9424 9126 9480
rect 9182 9424 65154 9480
rect 65210 9424 66166 9480
rect 66222 9424 66227 9480
rect 9121 9422 66227 9424
rect 9121 9419 9187 9422
rect 65149 9419 65215 9422
rect 66161 9419 66227 9422
rect 67398 9420 67404 9484
rect 67468 9482 67474 9484
rect 79041 9482 79107 9485
rect 67468 9480 79107 9482
rect 67468 9424 79046 9480
rect 79102 9424 79107 9480
rect 67468 9422 79107 9424
rect 67468 9420 67474 9422
rect 79041 9419 79107 9422
rect 79225 9482 79291 9485
rect 109534 9482 109540 9484
rect 79225 9480 109540 9482
rect 79225 9424 79230 9480
rect 79286 9424 109540 9480
rect 79225 9422 109540 9424
rect 79225 9419 79291 9422
rect 109534 9420 109540 9422
rect 109604 9420 109610 9484
rect 233734 9420 233740 9484
rect 233804 9482 233810 9484
rect 238710 9482 238770 9558
rect 233804 9422 238770 9482
rect 248137 9482 248203 9485
rect 248270 9482 248276 9484
rect 248137 9480 248276 9482
rect 248137 9424 248142 9480
rect 248198 9424 248276 9480
rect 248137 9422 248276 9424
rect 233804 9420 233810 9422
rect 248137 9419 248203 9422
rect 248270 9420 248276 9422
rect 248340 9420 248346 9484
rect 253890 9482 253950 9558
rect 272057 9616 273227 9618
rect 272057 9560 272062 9616
rect 272118 9560 273166 9616
rect 273222 9560 273227 9616
rect 272057 9558 273227 9560
rect 272057 9555 272123 9558
rect 273161 9555 273227 9558
rect 276606 9556 276612 9620
rect 276676 9618 276682 9620
rect 277761 9618 277827 9621
rect 276676 9616 277827 9618
rect 276676 9560 277766 9616
rect 277822 9560 277827 9616
rect 276676 9558 277827 9560
rect 276676 9556 276682 9558
rect 277761 9555 277827 9558
rect 273437 9482 273503 9485
rect 253890 9480 273503 9482
rect 253890 9424 273442 9480
rect 273498 9424 273503 9480
rect 253890 9422 273503 9424
rect 273437 9419 273503 9422
rect 35525 9346 35591 9349
rect 46054 9346 46060 9348
rect 35525 9344 46060 9346
rect 35525 9288 35530 9344
rect 35586 9288 46060 9344
rect 35525 9286 46060 9288
rect 35525 9283 35591 9286
rect 46054 9284 46060 9286
rect 46124 9284 46130 9348
rect 50286 9284 50292 9348
rect 50356 9346 50362 9348
rect 77937 9346 78003 9349
rect 50356 9344 78003 9346
rect 50356 9288 77942 9344
rect 77998 9288 78003 9344
rect 50356 9286 78003 9288
rect 50356 9284 50362 9286
rect 77937 9283 78003 9286
rect 78857 9346 78923 9349
rect 86166 9346 86172 9348
rect 78857 9344 86172 9346
rect 78857 9288 78862 9344
rect 78918 9288 86172 9344
rect 78857 9286 86172 9288
rect 78857 9283 78923 9286
rect 86166 9284 86172 9286
rect 86236 9284 86242 9348
rect 147070 9284 147076 9348
rect 147140 9346 147146 9348
rect 270861 9346 270927 9349
rect 273805 9346 273871 9349
rect 147140 9344 270927 9346
rect 147140 9288 270866 9344
rect 270922 9288 270927 9344
rect 147140 9286 270927 9288
rect 147140 9284 147146 9286
rect 270861 9283 270927 9286
rect 273210 9344 273871 9346
rect 273210 9288 273810 9344
rect 273866 9288 273871 9344
rect 273210 9286 273871 9288
rect 66161 9210 66227 9213
rect 222326 9210 222332 9212
rect 66161 9208 222332 9210
rect 66161 9152 66166 9208
rect 66222 9152 222332 9208
rect 66161 9150 222332 9152
rect 66161 9147 66227 9150
rect 222326 9148 222332 9150
rect 222396 9148 222402 9212
rect 230974 9148 230980 9212
rect 231044 9210 231050 9212
rect 240041 9210 240107 9213
rect 268326 9210 268332 9212
rect 231044 9208 240107 9210
rect 231044 9152 240046 9208
rect 240102 9152 240107 9208
rect 231044 9150 240107 9152
rect 231044 9148 231050 9150
rect 240041 9147 240107 9150
rect 248370 9150 268332 9210
rect 35014 9012 35020 9076
rect 35084 9074 35090 9076
rect 148041 9074 148107 9077
rect 35084 9072 148107 9074
rect 35084 9016 148046 9072
rect 148102 9016 148107 9072
rect 35084 9014 148107 9016
rect 35084 9012 35090 9014
rect 148041 9011 148107 9014
rect 239857 9074 239923 9077
rect 248370 9074 248430 9150
rect 268326 9148 268332 9150
rect 268396 9148 268402 9212
rect 270677 9210 270743 9213
rect 273210 9210 273270 9286
rect 273805 9283 273871 9286
rect 270677 9208 273270 9210
rect 270677 9152 270682 9208
rect 270738 9152 273270 9208
rect 270677 9150 273270 9152
rect 270677 9147 270743 9150
rect 239857 9072 248430 9074
rect 239857 9016 239862 9072
rect 239918 9016 248430 9072
rect 239857 9014 248430 9016
rect 272149 9074 272215 9077
rect 278129 9074 278195 9077
rect 272149 9072 278195 9074
rect 272149 9016 272154 9072
rect 272210 9016 278134 9072
rect 278190 9016 278195 9072
rect 272149 9014 278195 9016
rect 239857 9011 239923 9014
rect 272149 9011 272215 9014
rect 278129 9011 278195 9014
rect 77109 8938 77175 8941
rect 81934 8938 81940 8940
rect 77109 8936 81940 8938
rect -960 8802 480 8892
rect 77109 8880 77114 8936
rect 77170 8880 81940 8936
rect 77109 8878 81940 8880
rect 77109 8875 77175 8878
rect 81934 8876 81940 8878
rect 82004 8876 82010 8940
rect 88425 8938 88491 8941
rect 145782 8938 145788 8940
rect 88425 8936 145788 8938
rect 88425 8880 88430 8936
rect 88486 8880 145788 8936
rect 88425 8878 145788 8880
rect 88425 8875 88491 8878
rect 145782 8876 145788 8878
rect 145852 8876 145858 8940
rect 152549 8938 152615 8941
rect 207422 8938 207428 8940
rect 152549 8936 207428 8938
rect 152549 8880 152554 8936
rect 152610 8880 207428 8936
rect 152549 8878 207428 8880
rect 152549 8875 152615 8878
rect 207422 8876 207428 8878
rect 207492 8876 207498 8940
rect 270953 8938 271019 8941
rect 277577 8938 277643 8941
rect 270953 8936 277643 8938
rect 270953 8880 270958 8936
rect 271014 8880 277582 8936
rect 277638 8880 277643 8936
rect 270953 8878 277643 8880
rect 270953 8875 271019 8878
rect 277577 8875 277643 8878
rect 2773 8802 2839 8805
rect -960 8800 2839 8802
rect -960 8744 2778 8800
rect 2834 8744 2839 8800
rect -960 8742 2839 8744
rect -960 8652 480 8742
rect 2773 8739 2839 8742
rect 88609 8802 88675 8805
rect 125726 8802 125732 8804
rect 88609 8800 125732 8802
rect 88609 8744 88614 8800
rect 88670 8744 125732 8800
rect 88609 8742 125732 8744
rect 88609 8739 88675 8742
rect 125726 8740 125732 8742
rect 125796 8740 125802 8804
rect 196566 8740 196572 8804
rect 196636 8802 196642 8804
rect 244273 8802 244339 8805
rect 196636 8800 244339 8802
rect 196636 8744 244278 8800
rect 244334 8744 244339 8800
rect 196636 8742 244339 8744
rect 196636 8740 196642 8742
rect 244273 8739 244339 8742
rect 495433 8802 495499 8805
rect 499520 8802 500960 8892
rect 495433 8800 500960 8802
rect 495433 8744 495438 8800
rect 495494 8744 500960 8800
rect 495433 8742 500960 8744
rect 495433 8739 495499 8742
rect 3325 8666 3391 8669
rect 239857 8666 239923 8669
rect 3325 8664 239923 8666
rect 3325 8608 3330 8664
rect 3386 8608 239862 8664
rect 239918 8608 239923 8664
rect 499520 8652 500960 8742
rect 3325 8606 239923 8608
rect 3325 8603 3391 8606
rect 239857 8603 239923 8606
rect 88333 8530 88399 8533
rect 289670 8530 289676 8532
rect 88333 8528 289676 8530
rect 88333 8472 88338 8528
rect 88394 8472 289676 8528
rect 88333 8470 289676 8472
rect 88333 8467 88399 8470
rect 289670 8468 289676 8470
rect 289740 8468 289746 8532
rect 76414 8332 76420 8396
rect 76484 8394 76490 8396
rect 272333 8394 272399 8397
rect 76484 8392 272399 8394
rect 76484 8336 272338 8392
rect 272394 8336 272399 8392
rect 76484 8334 272399 8336
rect 76484 8332 76490 8334
rect 272333 8331 272399 8334
rect 76281 8258 76347 8261
rect 84326 8258 84332 8260
rect 76281 8256 84332 8258
rect 76281 8200 76286 8256
rect 76342 8200 84332 8256
rect 76281 8198 84332 8200
rect 76281 8195 76347 8198
rect 84326 8196 84332 8198
rect 84396 8196 84402 8260
rect 43161 8122 43227 8125
rect 53046 8122 53052 8124
rect 43161 8120 53052 8122
rect 43161 8064 43166 8120
rect 43222 8064 53052 8120
rect 43161 8062 53052 8064
rect 43161 8059 43227 8062
rect 53046 8060 53052 8062
rect 53116 8060 53122 8124
rect 57094 8060 57100 8124
rect 57164 8122 57170 8124
rect 109401 8122 109467 8125
rect 57164 8120 109467 8122
rect 57164 8064 109406 8120
rect 109462 8064 109467 8120
rect 57164 8062 109467 8064
rect 57164 8060 57170 8062
rect 109401 8059 109467 8062
rect 127566 8060 127572 8124
rect 127636 8122 127642 8124
rect 169017 8122 169083 8125
rect 127636 8120 169083 8122
rect 127636 8064 169022 8120
rect 169078 8064 169083 8120
rect 127636 8062 169083 8064
rect 127636 8060 127642 8062
rect 169017 8059 169083 8062
rect 3417 7986 3483 7989
rect 82905 7986 82971 7989
rect 3417 7984 82971 7986
rect 3417 7928 3422 7984
rect 3478 7928 82910 7984
rect 82966 7928 82971 7984
rect 3417 7926 82971 7928
rect 3417 7923 3483 7926
rect 82905 7923 82971 7926
rect 96153 7986 96219 7989
rect 112294 7986 112300 7988
rect 96153 7984 112300 7986
rect 96153 7928 96158 7984
rect 96214 7928 112300 7984
rect 96153 7926 112300 7928
rect 96153 7923 96219 7926
rect 112294 7924 112300 7926
rect 112364 7924 112370 7988
rect 116025 7986 116091 7989
rect 139894 7986 139900 7988
rect 116025 7984 139900 7986
rect 116025 7928 116030 7984
rect 116086 7928 139900 7984
rect 116025 7926 139900 7928
rect 116025 7923 116091 7926
rect 139894 7924 139900 7926
rect 139964 7924 139970 7988
rect 102777 7850 102843 7853
rect 180926 7850 180932 7852
rect 102777 7848 180932 7850
rect 102777 7792 102782 7848
rect 102838 7792 180932 7848
rect 102777 7790 180932 7792
rect 102777 7787 102843 7790
rect 180926 7788 180932 7790
rect 180996 7788 181002 7852
rect -960 4300 480 4540
rect 102869 4042 102935 4045
rect 104014 4042 104020 4044
rect 102869 4040 104020 4042
rect 102869 3984 102874 4040
rect 102930 3984 104020 4040
rect 102869 3982 104020 3984
rect 102869 3979 102935 3982
rect 104014 3980 104020 3982
rect 104084 3980 104090 4044
rect 123334 3980 123340 4044
rect 123404 4042 123410 4044
rect 178677 4042 178743 4045
rect 123404 4040 178743 4042
rect 123404 3984 178682 4040
rect 178738 3984 178743 4040
rect 123404 3982 178743 3984
rect 123404 3980 123410 3982
rect 178677 3979 178743 3982
rect 263358 3980 263364 4044
rect 263428 4042 263434 4044
rect 263501 4042 263567 4045
rect 263428 4040 263567 4042
rect 263428 3984 263506 4040
rect 263562 3984 263567 4040
rect 499520 4028 500960 4268
rect 263428 3982 263567 3984
rect 263428 3980 263434 3982
rect 263501 3979 263567 3982
rect 88190 3844 88196 3908
rect 88260 3906 88266 3908
rect 151445 3906 151511 3909
rect 88260 3904 151511 3906
rect 88260 3848 151450 3904
rect 151506 3848 151511 3904
rect 88260 3846 151511 3848
rect 88260 3844 88266 3846
rect 151445 3843 151511 3846
rect 98862 3708 98868 3772
rect 98932 3770 98938 3772
rect 100109 3770 100175 3773
rect 98932 3768 100175 3770
rect 98932 3712 100114 3768
rect 100170 3712 100175 3768
rect 98932 3710 100175 3712
rect 98932 3708 98938 3710
rect 100109 3707 100175 3710
rect 105997 3770 106063 3773
rect 108430 3770 108436 3772
rect 105997 3768 108436 3770
rect 105997 3712 106002 3768
rect 106058 3712 108436 3768
rect 105997 3710 108436 3712
rect 105997 3707 106063 3710
rect 108430 3708 108436 3710
rect 108500 3708 108506 3772
rect 124029 3770 124095 3773
rect 190310 3770 190316 3772
rect 124029 3768 190316 3770
rect 124029 3712 124034 3768
rect 124090 3712 190316 3768
rect 124029 3710 190316 3712
rect 124029 3707 124095 3710
rect 190310 3708 190316 3710
rect 190380 3708 190386 3772
rect 211981 3770 212047 3773
rect 212390 3770 212396 3772
rect 211981 3768 212396 3770
rect 211981 3712 211986 3768
rect 212042 3712 212396 3768
rect 211981 3710 212396 3712
rect 211981 3707 212047 3710
rect 212390 3708 212396 3710
rect 212460 3708 212466 3772
rect 217174 3708 217180 3772
rect 217244 3770 217250 3772
rect 266445 3770 266511 3773
rect 217244 3768 266511 3770
rect 217244 3712 266450 3768
rect 266506 3712 266511 3768
rect 217244 3710 266511 3712
rect 217244 3708 217250 3710
rect 266445 3707 266511 3710
rect 80646 3572 80652 3636
rect 80716 3634 80722 3636
rect 175549 3634 175615 3637
rect 80716 3632 175615 3634
rect 80716 3576 175554 3632
rect 175610 3576 175615 3632
rect 80716 3574 175615 3576
rect 80716 3572 80722 3574
rect 175549 3571 175615 3574
rect 190494 3572 190500 3636
rect 190564 3634 190570 3636
rect 242157 3634 242223 3637
rect 190564 3632 242223 3634
rect 190564 3576 242162 3632
rect 242218 3576 242223 3632
rect 190564 3574 242223 3576
rect 190564 3572 190570 3574
rect 242157 3571 242223 3574
rect 281533 3634 281599 3637
rect 375373 3634 375439 3637
rect 281533 3632 375439 3634
rect 281533 3576 281538 3632
rect 281594 3576 375378 3632
rect 375434 3576 375439 3632
rect 281533 3574 375439 3576
rect 281533 3571 281599 3574
rect 375373 3571 375439 3574
rect 36261 3498 36327 3501
rect 37774 3498 37780 3500
rect 36261 3496 37780 3498
rect 36261 3440 36266 3496
rect 36322 3440 37780 3496
rect 36261 3438 37780 3440
rect 36261 3435 36327 3438
rect 37774 3436 37780 3438
rect 37844 3436 37850 3500
rect 51349 3498 51415 3501
rect 52310 3498 52316 3500
rect 51349 3496 52316 3498
rect 51349 3440 51354 3496
rect 51410 3440 52316 3496
rect 51349 3438 52316 3440
rect 51349 3435 51415 3438
rect 52310 3436 52316 3438
rect 52380 3436 52386 3500
rect 72693 3498 72759 3501
rect 72918 3498 72924 3500
rect 72693 3496 72924 3498
rect 72693 3440 72698 3496
rect 72754 3440 72924 3496
rect 72693 3438 72924 3440
rect 72693 3435 72759 3438
rect 72918 3436 72924 3438
rect 72988 3436 72994 3500
rect 99414 3436 99420 3500
rect 99484 3498 99490 3500
rect 99925 3498 99991 3501
rect 99484 3496 99991 3498
rect 99484 3440 99930 3496
rect 99986 3440 99991 3496
rect 99484 3438 99991 3440
rect 99484 3436 99490 3438
rect 99925 3435 99991 3438
rect 100109 3498 100175 3501
rect 220997 3498 221063 3501
rect 100109 3496 221063 3498
rect 100109 3440 100114 3496
rect 100170 3440 221002 3496
rect 221058 3440 221063 3496
rect 100109 3438 221063 3440
rect 100109 3435 100175 3438
rect 220997 3435 221063 3438
rect 243486 3436 243492 3500
rect 243556 3498 243562 3500
rect 251357 3498 251423 3501
rect 243556 3496 251423 3498
rect 243556 3440 251362 3496
rect 251418 3440 251423 3496
rect 243556 3438 251423 3440
rect 243556 3436 243562 3438
rect 251357 3435 251423 3438
rect 313917 3498 313983 3501
rect 478413 3498 478479 3501
rect 313917 3496 478479 3498
rect 313917 3440 313922 3496
rect 313978 3440 478418 3496
rect 478474 3440 478479 3496
rect 313917 3438 478479 3440
rect 313917 3435 313983 3438
rect 478413 3435 478479 3438
rect 11973 3362 12039 3365
rect 415485 3362 415551 3365
rect 11973 3360 415551 3362
rect 11973 3304 11978 3360
rect 12034 3304 415490 3360
rect 415546 3304 415551 3360
rect 11973 3302 415551 3304
rect 11973 3299 12039 3302
rect 415485 3299 415551 3302
rect 138790 3164 138796 3228
rect 138860 3226 138866 3228
rect 169477 3226 169543 3229
rect 138860 3224 169543 3226
rect 138860 3168 169482 3224
rect 169538 3168 169543 3224
rect 138860 3166 169543 3168
rect 138860 3164 138866 3166
rect 169477 3163 169543 3166
rect 119654 3028 119660 3092
rect 119724 3090 119730 3092
rect 142245 3090 142311 3093
rect 119724 3088 142311 3090
rect 119724 3032 142250 3088
rect 142306 3032 142311 3088
rect 119724 3030 142311 3032
rect 119724 3028 119730 3030
rect 142245 3027 142311 3030
<< via3 >>
rect 90772 616796 90836 616860
rect 232452 616796 232516 616860
rect 234660 616796 234724 616860
rect 246252 616796 246316 616860
rect 295380 616856 295444 616860
rect 295380 616800 295394 616856
rect 295394 616800 295444 616856
rect 295380 616796 295444 616800
rect 184060 616252 184124 616316
rect 105492 616116 105556 616180
rect 258028 615572 258092 615636
rect 283420 610056 283484 610060
rect 283420 610000 283434 610056
rect 283434 610000 283484 610056
rect 283420 609996 283484 610000
rect 228588 606052 228652 606116
rect 50292 598980 50356 599044
rect 70900 596396 70964 596460
rect 205956 596320 206020 596324
rect 205956 596264 205970 596320
rect 205970 596264 206020 596320
rect 205956 596260 206020 596264
rect 201540 583808 201604 583812
rect 201540 583752 201554 583808
rect 201554 583752 201604 583808
rect 201540 583748 201604 583752
rect 111012 566068 111076 566132
rect 76420 565796 76484 565860
rect 268332 553480 268396 553484
rect 268332 553424 268346 553480
rect 268346 553424 268396 553480
rect 268332 553420 268396 553424
rect 276612 553420 276676 553484
rect 157564 543764 157628 543828
rect 123340 541648 123404 541652
rect 123340 541592 123354 541648
rect 123354 541592 123404 541648
rect 123340 541588 123404 541592
rect 128860 541452 128924 541516
rect 159220 539548 159284 539612
rect 117084 525268 117148 525332
rect 139900 525132 139964 525196
rect 96476 518740 96540 518804
rect 112300 518604 112364 518668
rect 190316 499624 190380 499628
rect 190316 499568 190366 499624
rect 190366 499568 190380 499624
rect 190316 499564 190380 499568
rect 220860 498068 220924 498132
rect 57100 493036 57164 493100
rect 32444 492688 32508 492692
rect 32444 492632 32458 492688
rect 32458 492632 32508 492688
rect 32444 492628 32508 492632
rect 145420 473452 145484 473516
rect 200620 470596 200684 470660
rect 146892 446932 146956 446996
rect 155172 442988 155236 443052
rect 263732 436112 263796 436116
rect 263732 436056 263746 436112
rect 263746 436056 263796 436112
rect 263732 436052 263796 436056
rect 34284 434964 34348 435028
rect 48084 434752 48148 434756
rect 48084 434696 48098 434752
rect 48098 434696 48148 434752
rect 48084 434692 48148 434696
rect 86172 433332 86236 433396
rect 36492 432108 36556 432172
rect 282684 432032 282748 432036
rect 282684 431976 282734 432032
rect 282734 431976 282748 432032
rect 282684 431972 282748 431976
rect 119660 414080 119724 414084
rect 119660 414024 119674 414080
rect 119674 414024 119724 414080
rect 119660 414020 119724 414024
rect 48820 410484 48884 410548
rect 55444 409940 55508 410004
rect 67404 400616 67468 400620
rect 67404 400560 67418 400616
rect 67418 400560 67468 400616
rect 67404 400556 67468 400560
rect 69612 400284 69676 400348
rect 132724 384236 132788 384300
rect 103652 384100 103716 384164
rect 88932 383964 88996 384028
rect 37780 383828 37844 383892
rect 38884 380972 38948 381036
rect 72924 380428 72988 380492
rect 233740 371784 233804 371788
rect 233740 371728 233754 371784
rect 233754 371728 233804 371784
rect 233740 371724 233804 371728
rect 217180 369820 217244 369884
rect 143212 365332 143276 365396
rect 196572 362476 196636 362540
rect 99420 356492 99484 356556
rect 117820 353364 117884 353428
rect 223620 337588 223684 337652
rect 230980 337376 231044 337380
rect 230980 337320 231030 337376
rect 231030 337320 231044 337376
rect 230980 337316 231044 337320
rect 38884 333296 38948 333300
rect 38884 333240 38898 333296
rect 38898 333240 38948 333296
rect 38884 333236 38948 333240
rect 263364 324940 263428 325004
rect 149652 306988 149716 307052
rect 261156 300928 261220 300932
rect 261156 300872 261170 300928
rect 261170 300872 261220 300928
rect 261156 300868 261220 300872
rect 113772 295564 113836 295628
rect 46060 288084 46124 288148
rect 108252 288084 108316 288148
rect 109540 286996 109604 287060
rect 274036 285696 274100 285700
rect 274036 285640 274050 285696
rect 274050 285640 274100 285696
rect 274036 285636 274100 285640
rect 191052 273804 191116 273868
rect 248276 273864 248340 273868
rect 248276 273808 248290 273864
rect 248290 273808 248340 273864
rect 248276 273804 248340 273808
rect 216076 267820 216140 267884
rect 103468 266928 103532 266932
rect 103468 266872 103482 266928
rect 103482 266872 103532 266928
rect 103468 266868 103532 266872
rect 98868 263604 98932 263668
rect 207428 262440 207492 262444
rect 207428 262384 207442 262440
rect 207442 262384 207492 262440
rect 207428 262380 207492 262384
rect 130332 261156 130396 261220
rect 125732 260884 125796 260948
rect 131620 260944 131684 260948
rect 131620 260888 131634 260944
rect 131634 260888 131684 260944
rect 131620 260884 131684 260888
rect 103284 259116 103348 259180
rect 180932 258572 180996 258636
rect 40540 254764 40604 254828
rect 219204 254688 219268 254692
rect 219204 254632 219254 254688
rect 219254 254632 219268 254688
rect 219204 254628 219268 254632
rect 303292 249868 303356 249932
rect 103468 248432 103532 248436
rect 103468 248376 103482 248432
rect 103482 248376 103532 248432
rect 103468 248372 103532 248376
rect 103652 238580 103716 238644
rect 62620 236132 62684 236196
rect 61516 236056 61580 236060
rect 61516 236000 61530 236056
rect 61530 236000 61580 236056
rect 61516 235996 61580 236000
rect 212396 232460 212460 232524
rect 188292 229740 188356 229804
rect 103468 229120 103532 229124
rect 103468 229064 103482 229120
rect 103482 229064 103532 229120
rect 103468 229060 103532 229064
rect 103468 228984 103532 228988
rect 103468 228928 103482 228984
rect 103482 228928 103532 228984
rect 103468 228924 103532 228928
rect 44036 228244 44100 228308
rect 53052 228108 53116 228172
rect 175780 228168 175844 228172
rect 175780 228112 175830 228168
rect 175830 228112 175844 228168
rect 175780 228108 175844 228112
rect 135668 227080 135732 227084
rect 135668 227024 135682 227080
rect 135682 227024 135732 227080
rect 135668 227020 135732 227024
rect 138612 226612 138676 226676
rect 103468 224904 103532 224908
rect 103468 224848 103482 224904
rect 103482 224848 103532 224904
rect 103468 224844 103532 224848
rect 63724 224436 63788 224500
rect 289676 223680 289740 223684
rect 289676 223624 289690 223680
rect 289690 223624 289740 223680
rect 289676 223620 289740 223624
rect 224724 222396 224788 222460
rect 59124 222260 59188 222324
rect 83964 222260 84028 222324
rect 204116 222260 204180 222324
rect 127572 220764 127636 220828
rect 209084 220824 209148 220828
rect 209084 220768 209098 220824
rect 209098 220768 209148 220824
rect 209084 220764 209148 220768
rect 124812 220628 124876 220692
rect 213132 220416 213196 220420
rect 213132 220360 213182 220416
rect 213182 220360 213196 220416
rect 213132 220356 213196 220360
rect 34468 219948 34532 220012
rect 42012 220008 42076 220012
rect 42012 219952 42062 220008
rect 42062 219952 42076 220008
rect 42012 219948 42076 219952
rect 51580 219948 51644 220012
rect 54340 219948 54404 220012
rect 68140 219948 68204 220012
rect 79548 219948 79612 220012
rect 94452 220008 94516 220012
rect 94452 219952 94502 220008
rect 94502 219952 94516 220008
rect 94452 219948 94516 219952
rect 101260 219948 101324 220012
rect 134380 219948 134444 220012
rect 153700 219948 153764 220012
rect 186820 219948 186884 220012
rect 193076 219948 193140 220012
rect 226932 220008 226996 220012
rect 226932 219952 226982 220008
rect 226982 219952 226996 220008
rect 226932 219948 226996 219952
rect 243492 219948 243556 220012
rect 253060 219948 253124 220012
rect 280660 219948 280724 220012
rect 77892 219812 77956 219876
rect 80652 219676 80716 219740
rect 240180 219736 240244 219740
rect 240180 219680 240194 219736
rect 240194 219680 240244 219736
rect 240180 219676 240244 219680
rect 162532 219540 162596 219604
rect 205036 219540 205100 219604
rect 87460 219404 87524 219468
rect 96660 219464 96724 219468
rect 96660 219408 96674 219464
rect 96674 219408 96724 219464
rect 96660 219404 96724 219408
rect 115060 219404 115124 219468
rect 162900 219404 162964 219468
rect 172468 219404 172532 219468
rect 173940 219464 174004 219468
rect 173940 219408 173990 219464
rect 173990 219408 174004 219464
rect 173940 219404 174004 219408
rect 184980 219404 185044 219468
rect 235948 219404 236012 219468
rect 273116 219404 273180 219468
rect 293172 219464 293236 219468
rect 293172 219408 293222 219464
rect 293222 219408 293236 219464
rect 293172 219404 293236 219408
rect 219388 219268 219452 219332
rect 210004 218588 210068 218652
rect 219020 121348 219084 121412
rect 219572 121348 219636 121412
rect 44036 120668 44100 120732
rect 96476 120728 96540 120732
rect 96476 120672 96490 120728
rect 96490 120672 96540 120728
rect 96476 120668 96540 120672
rect 103284 120668 103348 120732
rect 117084 120668 117148 120732
rect 34284 119988 34348 120052
rect 38884 119988 38948 120052
rect 55444 119988 55508 120052
rect 63724 120048 63788 120052
rect 63724 119992 63738 120048
rect 63738 119992 63788 120048
rect 63724 119988 63788 119992
rect 131620 119988 131684 120052
rect 258028 119988 258092 120052
rect 143212 119852 143276 119916
rect 162532 119912 162596 119916
rect 162532 119856 162546 119912
rect 162546 119856 162596 119912
rect 162532 119852 162596 119856
rect 200620 119852 200684 119916
rect 62620 119716 62684 119780
rect 61516 119580 61580 119644
rect 219204 119580 219268 119644
rect 216076 119504 216140 119508
rect 216076 119448 216090 119504
rect 216090 119448 216140 119504
rect 216076 119444 216140 119448
rect 40540 119308 40604 119372
rect 228588 119308 228652 119372
rect 263732 119308 263796 119372
rect 48084 119232 48148 119236
rect 48084 119176 48134 119232
rect 48134 119176 48148 119232
rect 48084 119172 48148 119176
rect 104020 119172 104084 119236
rect 36492 119036 36556 119100
rect 135668 119036 135732 119100
rect 145788 119036 145852 119100
rect 157564 119096 157628 119100
rect 157564 119040 157578 119096
rect 157578 119040 157628 119096
rect 157564 119036 157628 119040
rect 215892 119096 215956 119100
rect 215892 119040 215906 119096
rect 215906 119040 215956 119096
rect 215892 119036 215956 119040
rect 282684 118900 282748 118964
rect 35020 118764 35084 118828
rect 48820 118764 48884 118828
rect 147076 118764 147140 118828
rect 261340 118628 261404 118692
rect 234660 118492 234724 118556
rect 295380 118492 295444 118556
rect 32444 118356 32508 118420
rect 113772 118356 113836 118420
rect 253980 118356 254044 118420
rect 55812 118084 55876 118148
rect 79548 118220 79612 118284
rect 205036 118220 205100 118284
rect 223620 118220 223684 118284
rect 246252 118220 246316 118284
rect 84332 118084 84396 118148
rect 103284 118084 103348 118148
rect 141924 118084 141988 118148
rect 208900 118084 208964 118148
rect 269068 118084 269132 118148
rect 223620 117948 223684 118012
rect 249012 117948 249076 118012
rect 28764 117812 28828 117876
rect 121316 117812 121380 117876
rect 283420 117676 283484 117740
rect 293908 117676 293972 117740
rect 36492 117404 36556 117468
rect 49556 117404 49620 117468
rect 62620 117404 62684 117468
rect 82860 117404 82924 117468
rect 135852 117404 135916 117468
rect 149836 117404 149900 117468
rect 155356 117404 155420 117468
rect 161980 117404 162044 117468
rect 175964 117464 176028 117468
rect 175964 117408 175978 117464
rect 175978 117408 176028 117464
rect 175964 117404 176028 117408
rect 185164 117404 185228 117468
rect 188844 117404 188908 117468
rect 195100 117404 195164 117468
rect 202092 117404 202156 117468
rect 228220 117404 228284 117468
rect 235764 117404 235828 117468
rect 241652 117464 241716 117468
rect 241652 117408 241702 117464
rect 241702 117408 241716 117464
rect 241652 117404 241716 117408
rect 282132 117404 282196 117468
rect 287100 117268 287164 117332
rect 210004 115772 210068 115836
rect 70900 114412 70964 114476
rect 303292 113868 303356 113932
rect 186820 113052 186884 113116
rect 193076 113052 193140 113116
rect 219388 113052 219452 113116
rect 226932 113052 226996 113116
rect 273116 113052 273180 113116
rect 162900 112780 162964 112844
rect 172468 112780 172532 112844
rect 146892 112644 146956 112708
rect 225092 112644 225156 112708
rect 96660 112508 96724 112572
rect 201540 112508 201604 112572
rect 205956 112508 206020 112572
rect 149652 112372 149716 112436
rect 184980 112236 185044 112300
rect 52316 112100 52380 112164
rect 34468 111964 34532 112028
rect 42012 111964 42076 112028
rect 54340 111964 54404 112028
rect 59124 112100 59188 112164
rect 68140 112160 68204 112164
rect 68140 112104 68190 112160
rect 68190 112104 68204 112160
rect 68140 112100 68204 112104
rect 115060 112160 115124 112164
rect 115060 112104 115110 112160
rect 115110 112104 115124 112160
rect 115060 112100 115124 112104
rect 134380 112160 134444 112164
rect 134380 112104 134430 112160
rect 134430 112104 134444 112160
rect 134380 112100 134444 112104
rect 145420 112100 145484 112164
rect 153700 112100 153764 112164
rect 83964 111964 84028 112028
rect 87460 111964 87524 112028
rect 94452 111964 94516 112028
rect 101260 112024 101324 112028
rect 101260 111968 101310 112024
rect 101310 111968 101324 112024
rect 101260 111964 101324 111968
rect 108436 111964 108500 112028
rect 173940 111828 174004 111892
rect 204116 111828 204180 111892
rect 235948 111828 236012 111892
rect 240180 111828 240244 111892
rect 253060 111828 253124 111892
rect 280660 111828 280724 111892
rect 293172 111828 293236 111892
rect 159220 111692 159284 111756
rect 132724 111616 132788 111620
rect 132724 111560 132774 111616
rect 132774 111560 132788 111616
rect 132724 111556 132788 111560
rect 138612 111556 138676 111620
rect 130332 111420 130396 111484
rect 213132 111420 213196 111484
rect 128860 111284 128924 111348
rect 188292 111284 188356 111348
rect 111012 111148 111076 111212
rect 191052 111148 191116 111212
rect 232452 111148 232516 111212
rect 124812 111012 124876 111076
rect 274036 111012 274100 111076
rect 220860 110876 220924 110940
rect 51580 110740 51644 110804
rect 175780 110740 175844 110804
rect 90772 110604 90836 110668
rect 108252 110604 108316 110668
rect 138796 110468 138860 110532
rect 155172 110468 155236 110532
rect 182588 110528 182652 110532
rect 182588 110472 182638 110528
rect 182638 110472 182652 110528
rect 182588 110468 182652 110472
rect 190500 110528 190564 110532
rect 190500 110472 190514 110528
rect 190514 110472 190564 110528
rect 190500 110468 190564 110472
rect 209084 110468 209148 110532
rect 222332 110468 222396 110532
rect 273668 110528 273732 110532
rect 273668 110472 273682 110528
rect 273682 110472 273732 110528
rect 273668 110468 273732 110472
rect 88196 109440 88260 109444
rect 88196 109384 88210 109440
rect 88210 109384 88260 109440
rect 88196 109380 88260 109384
rect 293908 109108 293972 109172
rect 81940 108292 82004 108356
rect 182588 108292 182652 108356
rect 28764 10644 28828 10708
rect 49556 10644 49620 10708
rect 55812 10644 55876 10708
rect 62620 10644 62684 10708
rect 121316 10644 121380 10708
rect 155356 10644 155420 10708
rect 161980 10644 162044 10708
rect 175964 10704 176028 10708
rect 175964 10648 175978 10704
rect 175978 10648 176028 10704
rect 175964 10644 176028 10648
rect 185164 10644 185228 10708
rect 188844 10644 188908 10708
rect 195100 10644 195164 10708
rect 202092 10644 202156 10708
rect 208900 10704 208964 10708
rect 208900 10648 208914 10704
rect 208914 10648 208964 10704
rect 208900 10644 208964 10648
rect 228220 10644 228284 10708
rect 235764 10644 235828 10708
rect 249012 10644 249076 10708
rect 253980 10644 254044 10708
rect 261340 10644 261404 10708
rect 269068 10644 269132 10708
rect 273668 10644 273732 10708
rect 282132 10644 282196 10708
rect 287100 10644 287164 10708
rect 293908 10644 293972 10708
rect 215892 10236 215956 10300
rect 149836 10100 149900 10164
rect 241652 10160 241716 10164
rect 241652 10104 241702 10160
rect 241702 10104 241716 10160
rect 241652 10100 241716 10104
rect 36492 9888 36556 9892
rect 36492 9832 36542 9888
rect 36542 9832 36556 9888
rect 36492 9828 36556 9832
rect 82860 9888 82924 9892
rect 82860 9832 82910 9888
rect 82910 9832 82924 9888
rect 82860 9828 82924 9832
rect 135852 9888 135916 9892
rect 135852 9832 135902 9888
rect 135902 9832 135916 9888
rect 135852 9828 135916 9832
rect 142108 9828 142172 9892
rect 69612 9556 69676 9620
rect 77892 9616 77956 9620
rect 77892 9560 77906 9616
rect 77906 9560 77956 9616
rect 77892 9556 77956 9560
rect 88932 9556 88996 9620
rect 105492 9556 105556 9620
rect 117820 9556 117884 9620
rect 184060 9556 184124 9620
rect 67404 9420 67468 9484
rect 109540 9420 109604 9484
rect 233740 9420 233804 9484
rect 248276 9420 248340 9484
rect 276612 9556 276676 9620
rect 46060 9284 46124 9348
rect 50292 9284 50356 9348
rect 86172 9284 86236 9348
rect 147076 9284 147140 9348
rect 222332 9148 222396 9212
rect 230980 9148 231044 9212
rect 35020 9012 35084 9076
rect 268332 9148 268396 9212
rect 81940 8876 82004 8940
rect 145788 8876 145852 8940
rect 207428 8876 207492 8940
rect 125732 8740 125796 8804
rect 196572 8740 196636 8804
rect 289676 8468 289740 8532
rect 76420 8332 76484 8396
rect 84332 8196 84396 8260
rect 53052 8060 53116 8124
rect 57100 8060 57164 8124
rect 127572 8060 127636 8124
rect 112300 7924 112364 7988
rect 139900 7924 139964 7988
rect 180932 7788 180996 7852
rect 104020 3980 104084 4044
rect 123340 3980 123404 4044
rect 263364 3980 263428 4044
rect 88196 3844 88260 3908
rect 98868 3708 98932 3772
rect 108436 3708 108500 3772
rect 190316 3708 190380 3772
rect 212396 3708 212460 3772
rect 217180 3708 217244 3772
rect 80652 3572 80716 3636
rect 190500 3572 190564 3636
rect 37780 3436 37844 3500
rect 52316 3436 52380 3500
rect 72924 3436 72988 3500
rect 99420 3436 99484 3500
rect 243492 3436 243556 3500
rect 138796 3164 138860 3228
rect 119660 3028 119724 3092
<< metal4 >>
rect 90771 616860 90837 616861
rect 90771 616796 90772 616860
rect 90836 616796 90837 616860
rect 90771 616795 90837 616796
rect 232451 616860 232517 616861
rect 232451 616796 232452 616860
rect 232516 616796 232517 616860
rect 232451 616795 232517 616796
rect 234659 616860 234725 616861
rect 234659 616796 234660 616860
rect 234724 616796 234725 616860
rect 234659 616795 234725 616796
rect 246251 616860 246317 616861
rect 246251 616796 246252 616860
rect 246316 616796 246317 616860
rect 246251 616795 246317 616796
rect 295379 616860 295445 616861
rect 295379 616796 295380 616860
rect 295444 616796 295445 616860
rect 295379 616795 295445 616796
rect 50291 599044 50357 599045
rect 50291 598980 50292 599044
rect 50356 598980 50357 599044
rect 50291 598979 50357 598980
rect 32443 492692 32509 492693
rect 32443 492628 32444 492692
rect 32508 492628 32509 492692
rect 32443 492627 32509 492628
rect 32446 118421 32506 492627
rect 34283 435028 34349 435029
rect 34283 434964 34284 435028
rect 34348 434964 34349 435028
rect 34283 434963 34349 434964
rect 34286 120053 34346 434963
rect 48083 434756 48149 434757
rect 48083 434692 48084 434756
rect 48148 434692 48149 434756
rect 48083 434691 48149 434692
rect 36491 432172 36557 432173
rect 36491 432108 36492 432172
rect 36556 432108 36557 432172
rect 36491 432107 36557 432108
rect 34467 220012 34533 220013
rect 34467 219948 34468 220012
rect 34532 219948 34533 220012
rect 34467 219947 34533 219948
rect 34283 120052 34349 120053
rect 34283 119988 34284 120052
rect 34348 119988 34349 120052
rect 34283 119987 34349 119988
rect 32443 118420 32509 118421
rect 32443 118356 32444 118420
rect 32508 118356 32509 118420
rect 32443 118355 32509 118356
rect 28763 117876 28829 117877
rect 28763 117812 28764 117876
rect 28828 117812 28829 117876
rect 28763 117811 28829 117812
rect 28766 10709 28826 117811
rect 34470 112029 34530 219947
rect 36494 119101 36554 432107
rect 37779 383892 37845 383893
rect 37779 383828 37780 383892
rect 37844 383828 37845 383892
rect 37779 383827 37845 383828
rect 36491 119100 36557 119101
rect 36491 119036 36492 119100
rect 36556 119036 36557 119100
rect 36491 119035 36557 119036
rect 35019 118828 35085 118829
rect 35019 118764 35020 118828
rect 35084 118764 35085 118828
rect 35019 118763 35085 118764
rect 34467 112028 34533 112029
rect 34467 111964 34468 112028
rect 34532 111964 34533 112028
rect 34467 111963 34533 111964
rect 28763 10708 28829 10709
rect 28763 10644 28764 10708
rect 28828 10644 28829 10708
rect 28763 10643 28829 10644
rect 35022 9077 35082 118763
rect 36491 117468 36557 117469
rect 36491 117404 36492 117468
rect 36556 117404 36557 117468
rect 36491 117403 36557 117404
rect 36494 9893 36554 117403
rect 36491 9892 36557 9893
rect 36491 9828 36492 9892
rect 36556 9828 36557 9892
rect 36491 9827 36557 9828
rect 35019 9076 35085 9077
rect 35019 9012 35020 9076
rect 35084 9012 35085 9076
rect 35019 9011 35085 9012
rect 37782 3501 37842 383827
rect 38883 381036 38949 381037
rect 38883 380972 38884 381036
rect 38948 380972 38949 381036
rect 38883 380971 38949 380972
rect 38886 333301 38946 380971
rect 38883 333300 38949 333301
rect 38883 333236 38884 333300
rect 38948 333236 38949 333300
rect 38883 333235 38949 333236
rect 38886 120053 38946 333235
rect 46059 288148 46125 288149
rect 46059 288084 46060 288148
rect 46124 288084 46125 288148
rect 46059 288083 46125 288084
rect 40539 254828 40605 254829
rect 40539 254764 40540 254828
rect 40604 254764 40605 254828
rect 40539 254763 40605 254764
rect 38883 120052 38949 120053
rect 38883 119988 38884 120052
rect 38948 119988 38949 120052
rect 38883 119987 38949 119988
rect 40542 119373 40602 254763
rect 44035 228308 44101 228309
rect 44035 228244 44036 228308
rect 44100 228244 44101 228308
rect 44035 228243 44101 228244
rect 42011 220012 42077 220013
rect 42011 219948 42012 220012
rect 42076 219948 42077 220012
rect 42011 219947 42077 219948
rect 40539 119372 40605 119373
rect 40539 119308 40540 119372
rect 40604 119308 40605 119372
rect 40539 119307 40605 119308
rect 42014 112029 42074 219947
rect 44038 120733 44098 228243
rect 44035 120732 44101 120733
rect 44035 120668 44036 120732
rect 44100 120668 44101 120732
rect 44035 120667 44101 120668
rect 42011 112028 42077 112029
rect 42011 111964 42012 112028
rect 42076 111964 42077 112028
rect 42011 111963 42077 111964
rect 46062 9349 46122 288083
rect 48086 119237 48146 434691
rect 48819 410548 48885 410549
rect 48819 410484 48820 410548
rect 48884 410484 48885 410548
rect 48819 410483 48885 410484
rect 48083 119236 48149 119237
rect 48083 119172 48084 119236
rect 48148 119172 48149 119236
rect 48083 119171 48149 119172
rect 48822 118829 48882 410483
rect 48819 118828 48885 118829
rect 48819 118764 48820 118828
rect 48884 118764 48885 118828
rect 48819 118763 48885 118764
rect 49555 117468 49621 117469
rect 49555 117404 49556 117468
rect 49620 117404 49621 117468
rect 49555 117403 49621 117404
rect 49558 10709 49618 117403
rect 49555 10708 49621 10709
rect 49555 10644 49556 10708
rect 49620 10644 49621 10708
rect 49555 10643 49621 10644
rect 50294 9349 50354 598979
rect 70899 596460 70965 596461
rect 70899 596396 70900 596460
rect 70964 596396 70965 596460
rect 70899 596395 70965 596396
rect 57099 493100 57165 493101
rect 57099 493036 57100 493100
rect 57164 493036 57165 493100
rect 57099 493035 57165 493036
rect 55443 410004 55509 410005
rect 55443 409940 55444 410004
rect 55508 409940 55509 410004
rect 55443 409939 55509 409940
rect 53051 228172 53117 228173
rect 53051 228108 53052 228172
rect 53116 228108 53117 228172
rect 53051 228107 53117 228108
rect 51579 220012 51645 220013
rect 51579 219948 51580 220012
rect 51644 219948 51645 220012
rect 51579 219947 51645 219948
rect 51582 110805 51642 219947
rect 52315 112164 52381 112165
rect 52315 112100 52316 112164
rect 52380 112100 52381 112164
rect 52315 112099 52381 112100
rect 51579 110804 51645 110805
rect 51579 110740 51580 110804
rect 51644 110740 51645 110804
rect 51579 110739 51645 110740
rect 46059 9348 46125 9349
rect 46059 9284 46060 9348
rect 46124 9284 46125 9348
rect 46059 9283 46125 9284
rect 50291 9348 50357 9349
rect 50291 9284 50292 9348
rect 50356 9284 50357 9348
rect 50291 9283 50357 9284
rect 52318 3501 52378 112099
rect 53054 8125 53114 228107
rect 54339 220012 54405 220013
rect 54339 219948 54340 220012
rect 54404 219948 54405 220012
rect 54339 219947 54405 219948
rect 54342 112029 54402 219947
rect 55446 120053 55506 409939
rect 55443 120052 55509 120053
rect 55443 119988 55444 120052
rect 55508 119988 55509 120052
rect 55443 119987 55509 119988
rect 55811 118148 55877 118149
rect 55811 118084 55812 118148
rect 55876 118084 55877 118148
rect 55811 118083 55877 118084
rect 54339 112028 54405 112029
rect 54339 111964 54340 112028
rect 54404 111964 54405 112028
rect 54339 111963 54405 111964
rect 55814 10709 55874 118083
rect 55811 10708 55877 10709
rect 55811 10644 55812 10708
rect 55876 10644 55877 10708
rect 55811 10643 55877 10644
rect 57102 8125 57162 493035
rect 67403 400620 67469 400621
rect 67403 400556 67404 400620
rect 67468 400556 67469 400620
rect 67403 400555 67469 400556
rect 62619 236196 62685 236197
rect 62619 236132 62620 236196
rect 62684 236132 62685 236196
rect 62619 236131 62685 236132
rect 61515 236060 61581 236061
rect 61515 235996 61516 236060
rect 61580 235996 61581 236060
rect 61515 235995 61581 235996
rect 59123 222324 59189 222325
rect 59123 222260 59124 222324
rect 59188 222260 59189 222324
rect 59123 222259 59189 222260
rect 59126 112165 59186 222259
rect 61518 119645 61578 235995
rect 62622 119781 62682 236131
rect 63723 224500 63789 224501
rect 63723 224436 63724 224500
rect 63788 224436 63789 224500
rect 63723 224435 63789 224436
rect 63726 120053 63786 224435
rect 63723 120052 63789 120053
rect 63723 119988 63724 120052
rect 63788 119988 63789 120052
rect 63723 119987 63789 119988
rect 62619 119780 62685 119781
rect 62619 119716 62620 119780
rect 62684 119716 62685 119780
rect 62619 119715 62685 119716
rect 61515 119644 61581 119645
rect 61515 119580 61516 119644
rect 61580 119580 61581 119644
rect 61515 119579 61581 119580
rect 62619 117468 62685 117469
rect 62619 117404 62620 117468
rect 62684 117404 62685 117468
rect 62619 117403 62685 117404
rect 59123 112164 59189 112165
rect 59123 112100 59124 112164
rect 59188 112100 59189 112164
rect 59123 112099 59189 112100
rect 62622 10709 62682 117403
rect 62619 10708 62685 10709
rect 62619 10644 62620 10708
rect 62684 10644 62685 10708
rect 62619 10643 62685 10644
rect 67406 9485 67466 400555
rect 69611 400348 69677 400349
rect 69611 400284 69612 400348
rect 69676 400284 69677 400348
rect 69611 400283 69677 400284
rect 68139 220012 68205 220013
rect 68139 219948 68140 220012
rect 68204 219948 68205 220012
rect 68139 219947 68205 219948
rect 68142 112165 68202 219947
rect 68139 112164 68205 112165
rect 68139 112100 68140 112164
rect 68204 112100 68205 112164
rect 68139 112099 68205 112100
rect 69614 9621 69674 400283
rect 70902 114477 70962 596395
rect 76419 565860 76485 565861
rect 76419 565796 76420 565860
rect 76484 565796 76485 565860
rect 76419 565795 76485 565796
rect 72923 380492 72989 380493
rect 72923 380428 72924 380492
rect 72988 380428 72989 380492
rect 72923 380427 72989 380428
rect 70899 114476 70965 114477
rect 70899 114412 70900 114476
rect 70964 114412 70965 114476
rect 70899 114411 70965 114412
rect 69611 9620 69677 9621
rect 69611 9556 69612 9620
rect 69676 9556 69677 9620
rect 69611 9555 69677 9556
rect 67403 9484 67469 9485
rect 67403 9420 67404 9484
rect 67468 9420 67469 9484
rect 67403 9419 67469 9420
rect 53051 8124 53117 8125
rect 53051 8060 53052 8124
rect 53116 8060 53117 8124
rect 53051 8059 53117 8060
rect 57099 8124 57165 8125
rect 57099 8060 57100 8124
rect 57164 8060 57165 8124
rect 57099 8059 57165 8060
rect 72926 3501 72986 380427
rect 76422 8397 76482 565795
rect 86171 433396 86237 433397
rect 86171 433332 86172 433396
rect 86236 433332 86237 433396
rect 86171 433331 86237 433332
rect 83963 222324 84029 222325
rect 83963 222260 83964 222324
rect 84028 222260 84029 222324
rect 83963 222259 84029 222260
rect 79547 220012 79613 220013
rect 79547 219948 79548 220012
rect 79612 219948 79613 220012
rect 79547 219947 79613 219948
rect 77891 219876 77957 219877
rect 77891 219812 77892 219876
rect 77956 219812 77957 219876
rect 77891 219811 77957 219812
rect 77894 9621 77954 219811
rect 79550 118285 79610 219947
rect 80651 219740 80717 219741
rect 80651 219676 80652 219740
rect 80716 219676 80717 219740
rect 80651 219675 80717 219676
rect 79547 118284 79613 118285
rect 79547 118220 79548 118284
rect 79612 118220 79613 118284
rect 79547 118219 79613 118220
rect 77891 9620 77957 9621
rect 77891 9556 77892 9620
rect 77956 9556 77957 9620
rect 77891 9555 77957 9556
rect 76419 8396 76485 8397
rect 76419 8332 76420 8396
rect 76484 8332 76485 8396
rect 76419 8331 76485 8332
rect 80654 3637 80714 219675
rect 82859 117468 82925 117469
rect 82859 117404 82860 117468
rect 82924 117404 82925 117468
rect 82859 117403 82925 117404
rect 81939 108356 82005 108357
rect 81939 108292 81940 108356
rect 82004 108292 82005 108356
rect 81939 108291 82005 108292
rect 81942 8941 82002 108291
rect 82862 9893 82922 117403
rect 83966 112029 84026 222259
rect 84331 118148 84397 118149
rect 84331 118084 84332 118148
rect 84396 118084 84397 118148
rect 84331 118083 84397 118084
rect 83963 112028 84029 112029
rect 83963 111964 83964 112028
rect 84028 111964 84029 112028
rect 83963 111963 84029 111964
rect 82859 9892 82925 9893
rect 82859 9828 82860 9892
rect 82924 9828 82925 9892
rect 82859 9827 82925 9828
rect 81939 8940 82005 8941
rect 81939 8876 81940 8940
rect 82004 8876 82005 8940
rect 81939 8875 82005 8876
rect 84334 8261 84394 118083
rect 86174 9349 86234 433331
rect 88931 384028 88997 384029
rect 88931 383964 88932 384028
rect 88996 383964 88997 384028
rect 88931 383963 88997 383964
rect 87459 219468 87525 219469
rect 87459 219404 87460 219468
rect 87524 219404 87525 219468
rect 87459 219403 87525 219404
rect 87462 112029 87522 219403
rect 87459 112028 87525 112029
rect 87459 111964 87460 112028
rect 87524 111964 87525 112028
rect 87459 111963 87525 111964
rect 88195 109444 88261 109445
rect 88195 109380 88196 109444
rect 88260 109380 88261 109444
rect 88195 109379 88261 109380
rect 86171 9348 86237 9349
rect 86171 9284 86172 9348
rect 86236 9284 86237 9348
rect 86171 9283 86237 9284
rect 84331 8260 84397 8261
rect 84331 8196 84332 8260
rect 84396 8196 84397 8260
rect 84331 8195 84397 8196
rect 88198 3909 88258 109379
rect 88934 9621 88994 383963
rect 90774 110669 90834 616795
rect 184059 616316 184125 616317
rect 184059 616252 184060 616316
rect 184124 616252 184125 616316
rect 184059 616251 184125 616252
rect 105491 616180 105557 616181
rect 105491 616116 105492 616180
rect 105556 616116 105557 616180
rect 105491 616115 105557 616116
rect 96475 518804 96541 518805
rect 96475 518740 96476 518804
rect 96540 518740 96541 518804
rect 96475 518739 96541 518740
rect 94451 220012 94517 220013
rect 94451 219948 94452 220012
rect 94516 219948 94517 220012
rect 94451 219947 94517 219948
rect 94454 112029 94514 219947
rect 96478 120733 96538 518739
rect 103651 384164 103717 384165
rect 103651 384100 103652 384164
rect 103716 384100 103717 384164
rect 103651 384099 103717 384100
rect 103654 383670 103714 384099
rect 103286 383610 103714 383670
rect 99419 356556 99485 356557
rect 99419 356492 99420 356556
rect 99484 356492 99485 356556
rect 99419 356491 99485 356492
rect 98867 263668 98933 263669
rect 98867 263604 98868 263668
rect 98932 263604 98933 263668
rect 98867 263603 98933 263604
rect 96659 219468 96725 219469
rect 96659 219404 96660 219468
rect 96724 219404 96725 219468
rect 96659 219403 96725 219404
rect 96475 120732 96541 120733
rect 96475 120668 96476 120732
rect 96540 120668 96541 120732
rect 96475 120667 96541 120668
rect 96662 112573 96722 219403
rect 96659 112572 96725 112573
rect 96659 112508 96660 112572
rect 96724 112508 96725 112572
rect 96659 112507 96725 112508
rect 94451 112028 94517 112029
rect 94451 111964 94452 112028
rect 94516 111964 94517 112028
rect 94451 111963 94517 111964
rect 90771 110668 90837 110669
rect 90771 110604 90772 110668
rect 90836 110604 90837 110668
rect 90771 110603 90837 110604
rect 88931 9620 88997 9621
rect 88931 9556 88932 9620
rect 88996 9556 88997 9620
rect 88931 9555 88997 9556
rect 88195 3908 88261 3909
rect 88195 3844 88196 3908
rect 88260 3844 88261 3908
rect 88195 3843 88261 3844
rect 98870 3773 98930 263603
rect 98867 3772 98933 3773
rect 98867 3708 98868 3772
rect 98932 3708 98933 3772
rect 98867 3707 98933 3708
rect 80651 3636 80717 3637
rect 80651 3572 80652 3636
rect 80716 3572 80717 3636
rect 80651 3571 80717 3572
rect 99422 3501 99482 356491
rect 103286 266930 103346 383610
rect 103467 266932 103533 266933
rect 103467 266930 103468 266932
rect 103286 266870 103468 266930
rect 103467 266868 103468 266870
rect 103532 266868 103533 266932
rect 103467 266867 103533 266868
rect 103283 259180 103349 259181
rect 103283 259116 103284 259180
rect 103348 259116 103349 259180
rect 103283 259115 103349 259116
rect 103286 248430 103346 259115
rect 103102 248370 103346 248430
rect 103467 248436 103533 248437
rect 103467 248372 103468 248436
rect 103532 248372 103533 248436
rect 103467 248371 103533 248372
rect 103102 238770 103162 248370
rect 103470 247890 103530 248371
rect 103286 247830 103530 247890
rect 103286 239050 103346 247830
rect 103286 238990 103714 239050
rect 103102 238710 103346 238770
rect 103286 224970 103346 238710
rect 103654 238645 103714 238990
rect 103651 238644 103717 238645
rect 103651 238580 103652 238644
rect 103716 238580 103717 238644
rect 103651 238579 103717 238580
rect 103467 229124 103533 229125
rect 103467 229060 103468 229124
rect 103532 229060 103533 229124
rect 103467 229059 103533 229060
rect 103470 228989 103530 229059
rect 103467 228988 103533 228989
rect 103467 228924 103468 228988
rect 103532 228924 103533 228988
rect 103467 228923 103533 228924
rect 103102 224910 103346 224970
rect 103102 222210 103162 224910
rect 103467 224908 103533 224909
rect 103467 224844 103468 224908
rect 103532 224844 103533 224908
rect 103467 224843 103533 224844
rect 102918 222150 103162 222210
rect 101259 220012 101325 220013
rect 101259 219948 101260 220012
rect 101324 219948 101325 220012
rect 101259 219947 101325 219948
rect 101262 112029 101322 219947
rect 102918 212550 102978 222150
rect 102918 212490 103162 212550
rect 103102 122850 103162 212490
rect 103470 205650 103530 224843
rect 103286 205590 103530 205650
rect 103286 200130 103346 205590
rect 103286 200070 103530 200130
rect 103470 199610 103530 200070
rect 103286 199550 103530 199610
rect 103286 190770 103346 199550
rect 103286 190710 103530 190770
rect 103470 190470 103530 190710
rect 103286 190410 103530 190470
rect 103286 180810 103346 190410
rect 103286 180750 103530 180810
rect 103470 180570 103530 180750
rect 103286 180510 103530 180570
rect 103286 171730 103346 180510
rect 103286 171670 103714 171730
rect 103654 171150 103714 171670
rect 103286 171090 103714 171150
rect 103286 161490 103346 171090
rect 103286 161430 103714 161490
rect 103654 160850 103714 161430
rect 103286 160790 103714 160850
rect 103286 152010 103346 160790
rect 103286 151950 103530 152010
rect 103470 151830 103530 151950
rect 103286 151770 103530 151830
rect 103286 142170 103346 151770
rect 103286 142110 103530 142170
rect 103470 141810 103530 142110
rect 103286 141750 103530 141810
rect 103286 132970 103346 141750
rect 103286 132910 103530 132970
rect 103470 132510 103530 132910
rect 103286 132450 103530 132510
rect 103286 123450 103346 132450
rect 103286 123390 103714 123450
rect 103102 122790 103346 122850
rect 103286 120733 103346 122790
rect 103283 120732 103349 120733
rect 103283 120668 103284 120732
rect 103348 120668 103349 120732
rect 103283 120667 103349 120668
rect 103654 120050 103714 123390
rect 103286 119990 103714 120050
rect 103286 118149 103346 119990
rect 104019 119236 104085 119237
rect 104019 119172 104020 119236
rect 104084 119172 104085 119236
rect 104019 119171 104085 119172
rect 103283 118148 103349 118149
rect 103283 118084 103284 118148
rect 103348 118084 103349 118148
rect 103283 118083 103349 118084
rect 101259 112028 101325 112029
rect 101259 111964 101260 112028
rect 101324 111964 101325 112028
rect 101259 111963 101325 111964
rect 104022 4045 104082 119171
rect 105494 9621 105554 616115
rect 111011 566132 111077 566133
rect 111011 566068 111012 566132
rect 111076 566068 111077 566132
rect 111011 566067 111077 566068
rect 108251 288148 108317 288149
rect 108251 288084 108252 288148
rect 108316 288084 108317 288148
rect 108251 288083 108317 288084
rect 108254 110669 108314 288083
rect 109539 287060 109605 287061
rect 109539 286996 109540 287060
rect 109604 286996 109605 287060
rect 109539 286995 109605 286996
rect 108435 112028 108501 112029
rect 108435 111964 108436 112028
rect 108500 111964 108501 112028
rect 108435 111963 108501 111964
rect 108251 110668 108317 110669
rect 108251 110604 108252 110668
rect 108316 110604 108317 110668
rect 108251 110603 108317 110604
rect 105491 9620 105557 9621
rect 105491 9556 105492 9620
rect 105556 9556 105557 9620
rect 105491 9555 105557 9556
rect 104019 4044 104085 4045
rect 104019 3980 104020 4044
rect 104084 3980 104085 4044
rect 104019 3979 104085 3980
rect 108438 3773 108498 111963
rect 109542 9485 109602 286995
rect 111014 111213 111074 566067
rect 157563 543828 157629 543829
rect 157563 543764 157564 543828
rect 157628 543764 157629 543828
rect 157563 543763 157629 543764
rect 123339 541652 123405 541653
rect 123339 541588 123340 541652
rect 123404 541588 123405 541652
rect 123339 541587 123405 541588
rect 117083 525332 117149 525333
rect 117083 525268 117084 525332
rect 117148 525268 117149 525332
rect 117083 525267 117149 525268
rect 112299 518668 112365 518669
rect 112299 518604 112300 518668
rect 112364 518604 112365 518668
rect 112299 518603 112365 518604
rect 111011 111212 111077 111213
rect 111011 111148 111012 111212
rect 111076 111148 111077 111212
rect 111011 111147 111077 111148
rect 109539 9484 109605 9485
rect 109539 9420 109540 9484
rect 109604 9420 109605 9484
rect 109539 9419 109605 9420
rect 112302 7989 112362 518603
rect 113771 295628 113837 295629
rect 113771 295564 113772 295628
rect 113836 295564 113837 295628
rect 113771 295563 113837 295564
rect 113774 118421 113834 295563
rect 115059 219468 115125 219469
rect 115059 219404 115060 219468
rect 115124 219404 115125 219468
rect 115059 219403 115125 219404
rect 113771 118420 113837 118421
rect 113771 118356 113772 118420
rect 113836 118356 113837 118420
rect 113771 118355 113837 118356
rect 115062 112165 115122 219403
rect 117086 120733 117146 525267
rect 119659 414084 119725 414085
rect 119659 414020 119660 414084
rect 119724 414020 119725 414084
rect 119659 414019 119725 414020
rect 117819 353428 117885 353429
rect 117819 353364 117820 353428
rect 117884 353364 117885 353428
rect 117819 353363 117885 353364
rect 117083 120732 117149 120733
rect 117083 120668 117084 120732
rect 117148 120668 117149 120732
rect 117083 120667 117149 120668
rect 115059 112164 115125 112165
rect 115059 112100 115060 112164
rect 115124 112100 115125 112164
rect 115059 112099 115125 112100
rect 117822 9621 117882 353363
rect 117819 9620 117885 9621
rect 117819 9556 117820 9620
rect 117884 9556 117885 9620
rect 117819 9555 117885 9556
rect 112299 7988 112365 7989
rect 112299 7924 112300 7988
rect 112364 7924 112365 7988
rect 112299 7923 112365 7924
rect 108435 3772 108501 3773
rect 108435 3708 108436 3772
rect 108500 3708 108501 3772
rect 108435 3707 108501 3708
rect 37779 3500 37845 3501
rect 37779 3436 37780 3500
rect 37844 3436 37845 3500
rect 37779 3435 37845 3436
rect 52315 3500 52381 3501
rect 52315 3436 52316 3500
rect 52380 3436 52381 3500
rect 52315 3435 52381 3436
rect 72923 3500 72989 3501
rect 72923 3436 72924 3500
rect 72988 3436 72989 3500
rect 72923 3435 72989 3436
rect 99419 3500 99485 3501
rect 99419 3436 99420 3500
rect 99484 3436 99485 3500
rect 99419 3435 99485 3436
rect 119662 3093 119722 414019
rect 121315 117876 121381 117877
rect 121315 117812 121316 117876
rect 121380 117812 121381 117876
rect 121315 117811 121381 117812
rect 121318 10709 121378 117811
rect 121315 10708 121381 10709
rect 121315 10644 121316 10708
rect 121380 10644 121381 10708
rect 121315 10643 121381 10644
rect 123342 4045 123402 541587
rect 128859 541516 128925 541517
rect 128859 541452 128860 541516
rect 128924 541452 128925 541516
rect 128859 541451 128925 541452
rect 125731 260948 125797 260949
rect 125731 260884 125732 260948
rect 125796 260884 125797 260948
rect 125731 260883 125797 260884
rect 124811 220692 124877 220693
rect 124811 220628 124812 220692
rect 124876 220628 124877 220692
rect 124811 220627 124877 220628
rect 124814 111077 124874 220627
rect 124811 111076 124877 111077
rect 124811 111012 124812 111076
rect 124876 111012 124877 111076
rect 124811 111011 124877 111012
rect 125734 8805 125794 260883
rect 127571 220828 127637 220829
rect 127571 220764 127572 220828
rect 127636 220764 127637 220828
rect 127571 220763 127637 220764
rect 125731 8804 125797 8805
rect 125731 8740 125732 8804
rect 125796 8740 125797 8804
rect 125731 8739 125797 8740
rect 127574 8125 127634 220763
rect 128862 111349 128922 541451
rect 139899 525196 139965 525197
rect 139899 525132 139900 525196
rect 139964 525132 139965 525196
rect 139899 525131 139965 525132
rect 132723 384300 132789 384301
rect 132723 384236 132724 384300
rect 132788 384236 132789 384300
rect 132723 384235 132789 384236
rect 130331 261220 130397 261221
rect 130331 261156 130332 261220
rect 130396 261156 130397 261220
rect 130331 261155 130397 261156
rect 130334 111485 130394 261155
rect 131619 260948 131685 260949
rect 131619 260884 131620 260948
rect 131684 260884 131685 260948
rect 131619 260883 131685 260884
rect 131622 120053 131682 260883
rect 131619 120052 131685 120053
rect 131619 119988 131620 120052
rect 131684 119988 131685 120052
rect 131619 119987 131685 119988
rect 132726 111621 132786 384235
rect 135667 227084 135733 227085
rect 135667 227020 135668 227084
rect 135732 227020 135733 227084
rect 135667 227019 135733 227020
rect 134379 220012 134445 220013
rect 134379 219948 134380 220012
rect 134444 219948 134445 220012
rect 134379 219947 134445 219948
rect 134382 112165 134442 219947
rect 135670 119101 135730 227019
rect 138611 226676 138677 226677
rect 138611 226612 138612 226676
rect 138676 226612 138677 226676
rect 138611 226611 138677 226612
rect 135667 119100 135733 119101
rect 135667 119036 135668 119100
rect 135732 119036 135733 119100
rect 135667 119035 135733 119036
rect 135851 117468 135917 117469
rect 135851 117404 135852 117468
rect 135916 117404 135917 117468
rect 135851 117403 135917 117404
rect 134379 112164 134445 112165
rect 134379 112100 134380 112164
rect 134444 112100 134445 112164
rect 134379 112099 134445 112100
rect 132723 111620 132789 111621
rect 132723 111556 132724 111620
rect 132788 111556 132789 111620
rect 132723 111555 132789 111556
rect 130331 111484 130397 111485
rect 130331 111420 130332 111484
rect 130396 111420 130397 111484
rect 130331 111419 130397 111420
rect 128859 111348 128925 111349
rect 128859 111284 128860 111348
rect 128924 111284 128925 111348
rect 128859 111283 128925 111284
rect 135854 9893 135914 117403
rect 138614 111621 138674 226611
rect 138611 111620 138677 111621
rect 138611 111556 138612 111620
rect 138676 111556 138677 111620
rect 138611 111555 138677 111556
rect 138795 110532 138861 110533
rect 138795 110468 138796 110532
rect 138860 110468 138861 110532
rect 138795 110467 138861 110468
rect 135851 9892 135917 9893
rect 135851 9828 135852 9892
rect 135916 9828 135917 9892
rect 135851 9827 135917 9828
rect 127571 8124 127637 8125
rect 127571 8060 127572 8124
rect 127636 8060 127637 8124
rect 127571 8059 127637 8060
rect 123339 4044 123405 4045
rect 123339 3980 123340 4044
rect 123404 3980 123405 4044
rect 123339 3979 123405 3980
rect 138798 3229 138858 110467
rect 139902 7989 139962 525131
rect 145419 473516 145485 473517
rect 145419 473452 145420 473516
rect 145484 473452 145485 473516
rect 145419 473451 145485 473452
rect 143211 365396 143277 365397
rect 143211 365332 143212 365396
rect 143276 365332 143277 365396
rect 143211 365331 143277 365332
rect 143214 119917 143274 365331
rect 143211 119916 143277 119917
rect 143211 119852 143212 119916
rect 143276 119852 143277 119916
rect 143211 119851 143277 119852
rect 141923 118148 141989 118149
rect 141923 118084 141924 118148
rect 141988 118084 141989 118148
rect 141923 118083 141989 118084
rect 141926 9890 141986 118083
rect 145422 112165 145482 473451
rect 146891 446996 146957 446997
rect 146891 446932 146892 446996
rect 146956 446932 146957 446996
rect 146891 446931 146957 446932
rect 145787 119100 145853 119101
rect 145787 119036 145788 119100
rect 145852 119036 145853 119100
rect 145787 119035 145853 119036
rect 145419 112164 145485 112165
rect 145419 112100 145420 112164
rect 145484 112100 145485 112164
rect 145419 112099 145485 112100
rect 142107 9892 142173 9893
rect 142107 9890 142108 9892
rect 141926 9830 142108 9890
rect 142107 9828 142108 9830
rect 142172 9828 142173 9892
rect 142107 9827 142173 9828
rect 145790 8941 145850 119035
rect 146894 112709 146954 446931
rect 155171 443052 155237 443053
rect 155171 442988 155172 443052
rect 155236 442988 155237 443052
rect 155171 442987 155237 442988
rect 149651 307052 149717 307053
rect 149651 306988 149652 307052
rect 149716 306988 149717 307052
rect 149651 306987 149717 306988
rect 147075 118828 147141 118829
rect 147075 118764 147076 118828
rect 147140 118764 147141 118828
rect 147075 118763 147141 118764
rect 146891 112708 146957 112709
rect 146891 112644 146892 112708
rect 146956 112644 146957 112708
rect 146891 112643 146957 112644
rect 147078 9349 147138 118763
rect 149654 112437 149714 306987
rect 153699 220012 153765 220013
rect 153699 219948 153700 220012
rect 153764 219948 153765 220012
rect 153699 219947 153765 219948
rect 149835 117468 149901 117469
rect 149835 117404 149836 117468
rect 149900 117404 149901 117468
rect 149835 117403 149901 117404
rect 149651 112436 149717 112437
rect 149651 112372 149652 112436
rect 149716 112372 149717 112436
rect 149651 112371 149717 112372
rect 149838 10165 149898 117403
rect 153702 112165 153762 219947
rect 153699 112164 153765 112165
rect 153699 112100 153700 112164
rect 153764 112100 153765 112164
rect 153699 112099 153765 112100
rect 155174 110533 155234 442987
rect 157566 119101 157626 543763
rect 159219 539612 159285 539613
rect 159219 539548 159220 539612
rect 159284 539548 159285 539612
rect 159219 539547 159285 539548
rect 157563 119100 157629 119101
rect 157563 119036 157564 119100
rect 157628 119036 157629 119100
rect 157563 119035 157629 119036
rect 155355 117468 155421 117469
rect 155355 117404 155356 117468
rect 155420 117404 155421 117468
rect 155355 117403 155421 117404
rect 155171 110532 155237 110533
rect 155171 110468 155172 110532
rect 155236 110468 155237 110532
rect 155171 110467 155237 110468
rect 155358 10709 155418 117403
rect 159222 111757 159282 539547
rect 180931 258636 180997 258637
rect 180931 258572 180932 258636
rect 180996 258572 180997 258636
rect 180931 258571 180997 258572
rect 175779 228172 175845 228173
rect 175779 228108 175780 228172
rect 175844 228108 175845 228172
rect 175779 228107 175845 228108
rect 162531 219604 162597 219605
rect 162531 219540 162532 219604
rect 162596 219540 162597 219604
rect 162531 219539 162597 219540
rect 162534 119917 162594 219539
rect 162899 219468 162965 219469
rect 162899 219404 162900 219468
rect 162964 219404 162965 219468
rect 162899 219403 162965 219404
rect 172467 219468 172533 219469
rect 172467 219404 172468 219468
rect 172532 219404 172533 219468
rect 172467 219403 172533 219404
rect 173939 219468 174005 219469
rect 173939 219404 173940 219468
rect 174004 219404 174005 219468
rect 173939 219403 174005 219404
rect 162531 119916 162597 119917
rect 162531 119852 162532 119916
rect 162596 119852 162597 119916
rect 162531 119851 162597 119852
rect 161979 117468 162045 117469
rect 161979 117404 161980 117468
rect 162044 117404 162045 117468
rect 161979 117403 162045 117404
rect 159219 111756 159285 111757
rect 159219 111692 159220 111756
rect 159284 111692 159285 111756
rect 159219 111691 159285 111692
rect 161982 10709 162042 117403
rect 162902 112845 162962 219403
rect 172470 112845 172530 219403
rect 162899 112844 162965 112845
rect 162899 112780 162900 112844
rect 162964 112780 162965 112844
rect 162899 112779 162965 112780
rect 172467 112844 172533 112845
rect 172467 112780 172468 112844
rect 172532 112780 172533 112844
rect 172467 112779 172533 112780
rect 173942 111893 174002 219403
rect 173939 111892 174005 111893
rect 173939 111828 173940 111892
rect 174004 111828 174005 111892
rect 173939 111827 174005 111828
rect 175782 110805 175842 228107
rect 175963 117468 176029 117469
rect 175963 117404 175964 117468
rect 176028 117404 176029 117468
rect 175963 117403 176029 117404
rect 175779 110804 175845 110805
rect 175779 110740 175780 110804
rect 175844 110740 175845 110804
rect 175779 110739 175845 110740
rect 175966 10709 176026 117403
rect 155355 10708 155421 10709
rect 155355 10644 155356 10708
rect 155420 10644 155421 10708
rect 155355 10643 155421 10644
rect 161979 10708 162045 10709
rect 161979 10644 161980 10708
rect 162044 10644 162045 10708
rect 161979 10643 162045 10644
rect 175963 10708 176029 10709
rect 175963 10644 175964 10708
rect 176028 10644 176029 10708
rect 175963 10643 176029 10644
rect 149835 10164 149901 10165
rect 149835 10100 149836 10164
rect 149900 10100 149901 10164
rect 149835 10099 149901 10100
rect 147075 9348 147141 9349
rect 147075 9284 147076 9348
rect 147140 9284 147141 9348
rect 147075 9283 147141 9284
rect 145787 8940 145853 8941
rect 145787 8876 145788 8940
rect 145852 8876 145853 8940
rect 145787 8875 145853 8876
rect 139899 7988 139965 7989
rect 139899 7924 139900 7988
rect 139964 7924 139965 7988
rect 139899 7923 139965 7924
rect 180934 7853 180994 258571
rect 182587 110532 182653 110533
rect 182587 110468 182588 110532
rect 182652 110468 182653 110532
rect 182587 110467 182653 110468
rect 182590 108357 182650 110467
rect 182587 108356 182653 108357
rect 182587 108292 182588 108356
rect 182652 108292 182653 108356
rect 182587 108291 182653 108292
rect 184062 9621 184122 616251
rect 228587 606116 228653 606117
rect 228587 606052 228588 606116
rect 228652 606052 228653 606116
rect 228587 606051 228653 606052
rect 205955 596324 206021 596325
rect 205955 596260 205956 596324
rect 206020 596260 206021 596324
rect 205955 596259 206021 596260
rect 201539 583812 201605 583813
rect 201539 583748 201540 583812
rect 201604 583748 201605 583812
rect 201539 583747 201605 583748
rect 190315 499628 190381 499629
rect 190315 499564 190316 499628
rect 190380 499564 190381 499628
rect 190315 499563 190381 499564
rect 188291 229804 188357 229805
rect 188291 229740 188292 229804
rect 188356 229740 188357 229804
rect 188291 229739 188357 229740
rect 186819 220012 186885 220013
rect 186819 219948 186820 220012
rect 186884 219948 186885 220012
rect 186819 219947 186885 219948
rect 184979 219468 185045 219469
rect 184979 219404 184980 219468
rect 185044 219404 185045 219468
rect 184979 219403 185045 219404
rect 184982 112301 185042 219403
rect 185163 117468 185229 117469
rect 185163 117404 185164 117468
rect 185228 117404 185229 117468
rect 185163 117403 185229 117404
rect 184979 112300 185045 112301
rect 184979 112236 184980 112300
rect 185044 112236 185045 112300
rect 184979 112235 185045 112236
rect 185166 10709 185226 117403
rect 186822 113117 186882 219947
rect 186819 113116 186885 113117
rect 186819 113052 186820 113116
rect 186884 113052 186885 113116
rect 186819 113051 186885 113052
rect 188294 111349 188354 229739
rect 188843 117468 188909 117469
rect 188843 117404 188844 117468
rect 188908 117404 188909 117468
rect 188843 117403 188909 117404
rect 188291 111348 188357 111349
rect 188291 111284 188292 111348
rect 188356 111284 188357 111348
rect 188291 111283 188357 111284
rect 188846 10709 188906 117403
rect 185163 10708 185229 10709
rect 185163 10644 185164 10708
rect 185228 10644 185229 10708
rect 185163 10643 185229 10644
rect 188843 10708 188909 10709
rect 188843 10644 188844 10708
rect 188908 10644 188909 10708
rect 188843 10643 188909 10644
rect 184059 9620 184125 9621
rect 184059 9556 184060 9620
rect 184124 9556 184125 9620
rect 184059 9555 184125 9556
rect 180931 7852 180997 7853
rect 180931 7788 180932 7852
rect 180996 7788 180997 7852
rect 180931 7787 180997 7788
rect 190318 3773 190378 499563
rect 200619 470660 200685 470661
rect 200619 470596 200620 470660
rect 200684 470596 200685 470660
rect 200619 470595 200685 470596
rect 196571 362540 196637 362541
rect 196571 362476 196572 362540
rect 196636 362476 196637 362540
rect 196571 362475 196637 362476
rect 191051 273868 191117 273869
rect 191051 273804 191052 273868
rect 191116 273804 191117 273868
rect 191051 273803 191117 273804
rect 191054 111213 191114 273803
rect 193075 220012 193141 220013
rect 193075 219948 193076 220012
rect 193140 219948 193141 220012
rect 193075 219947 193141 219948
rect 193078 113117 193138 219947
rect 195099 117468 195165 117469
rect 195099 117404 195100 117468
rect 195164 117404 195165 117468
rect 195099 117403 195165 117404
rect 193075 113116 193141 113117
rect 193075 113052 193076 113116
rect 193140 113052 193141 113116
rect 193075 113051 193141 113052
rect 191051 111212 191117 111213
rect 191051 111148 191052 111212
rect 191116 111148 191117 111212
rect 191051 111147 191117 111148
rect 190499 110532 190565 110533
rect 190499 110468 190500 110532
rect 190564 110468 190565 110532
rect 190499 110467 190565 110468
rect 190315 3772 190381 3773
rect 190315 3708 190316 3772
rect 190380 3708 190381 3772
rect 190315 3707 190381 3708
rect 190502 3637 190562 110467
rect 195102 10709 195162 117403
rect 195099 10708 195165 10709
rect 195099 10644 195100 10708
rect 195164 10644 195165 10708
rect 195099 10643 195165 10644
rect 196574 8805 196634 362475
rect 200622 119917 200682 470595
rect 200619 119916 200685 119917
rect 200619 119852 200620 119916
rect 200684 119852 200685 119916
rect 200619 119851 200685 119852
rect 201542 112573 201602 583747
rect 204115 222324 204181 222325
rect 204115 222260 204116 222324
rect 204180 222260 204181 222324
rect 204115 222259 204181 222260
rect 202091 117468 202157 117469
rect 202091 117404 202092 117468
rect 202156 117404 202157 117468
rect 202091 117403 202157 117404
rect 201539 112572 201605 112573
rect 201539 112508 201540 112572
rect 201604 112508 201605 112572
rect 201539 112507 201605 112508
rect 202094 10709 202154 117403
rect 204118 111893 204178 222259
rect 205035 219604 205101 219605
rect 205035 219540 205036 219604
rect 205100 219540 205101 219604
rect 205035 219539 205101 219540
rect 205038 118285 205098 219539
rect 205035 118284 205101 118285
rect 205035 118220 205036 118284
rect 205100 118220 205101 118284
rect 205035 118219 205101 118220
rect 205958 112573 206018 596259
rect 220859 498132 220925 498133
rect 220859 498068 220860 498132
rect 220924 498068 220925 498132
rect 220859 498067 220925 498068
rect 217179 369884 217245 369885
rect 217179 369820 217180 369884
rect 217244 369820 217245 369884
rect 217179 369819 217245 369820
rect 216075 267884 216141 267885
rect 216075 267820 216076 267884
rect 216140 267820 216141 267884
rect 216075 267819 216141 267820
rect 207427 262444 207493 262445
rect 207427 262380 207428 262444
rect 207492 262380 207493 262444
rect 207427 262379 207493 262380
rect 205955 112572 206021 112573
rect 205955 112508 205956 112572
rect 206020 112508 206021 112572
rect 205955 112507 206021 112508
rect 204115 111892 204181 111893
rect 204115 111828 204116 111892
rect 204180 111828 204181 111892
rect 204115 111827 204181 111828
rect 202091 10708 202157 10709
rect 202091 10644 202092 10708
rect 202156 10644 202157 10708
rect 202091 10643 202157 10644
rect 207430 8941 207490 262379
rect 212395 232524 212461 232525
rect 212395 232460 212396 232524
rect 212460 232460 212461 232524
rect 212395 232459 212461 232460
rect 209083 220828 209149 220829
rect 209083 220764 209084 220828
rect 209148 220764 209149 220828
rect 209083 220763 209149 220764
rect 208899 118148 208965 118149
rect 208899 118084 208900 118148
rect 208964 118084 208965 118148
rect 208899 118083 208965 118084
rect 208902 10709 208962 118083
rect 209086 110533 209146 220763
rect 210003 218652 210069 218653
rect 210003 218588 210004 218652
rect 210068 218588 210069 218652
rect 210003 218587 210069 218588
rect 210006 115837 210066 218587
rect 210003 115836 210069 115837
rect 210003 115772 210004 115836
rect 210068 115772 210069 115836
rect 210003 115771 210069 115772
rect 209083 110532 209149 110533
rect 209083 110468 209084 110532
rect 209148 110468 209149 110532
rect 209083 110467 209149 110468
rect 208899 10708 208965 10709
rect 208899 10644 208900 10708
rect 208964 10644 208965 10708
rect 208899 10643 208965 10644
rect 207427 8940 207493 8941
rect 207427 8876 207428 8940
rect 207492 8876 207493 8940
rect 207427 8875 207493 8876
rect 196571 8804 196637 8805
rect 196571 8740 196572 8804
rect 196636 8740 196637 8804
rect 196571 8739 196637 8740
rect 212398 3773 212458 232459
rect 213131 220420 213197 220421
rect 213131 220356 213132 220420
rect 213196 220356 213197 220420
rect 213131 220355 213197 220356
rect 213134 111485 213194 220355
rect 216078 119509 216138 267819
rect 216075 119508 216141 119509
rect 216075 119444 216076 119508
rect 216140 119444 216141 119508
rect 216075 119443 216141 119444
rect 215891 119100 215957 119101
rect 215891 119036 215892 119100
rect 215956 119036 215957 119100
rect 215891 119035 215957 119036
rect 213131 111484 213197 111485
rect 213131 111420 213132 111484
rect 213196 111420 213197 111484
rect 213131 111419 213197 111420
rect 215894 10301 215954 119035
rect 215891 10300 215957 10301
rect 215891 10236 215892 10300
rect 215956 10236 215957 10300
rect 215891 10235 215957 10236
rect 217182 3773 217242 369819
rect 219203 254692 219269 254693
rect 219203 254628 219204 254692
rect 219268 254628 219269 254692
rect 219203 254627 219269 254628
rect 219206 224970 219266 254627
rect 219022 224910 219266 224970
rect 219022 222210 219082 224910
rect 219022 222150 219266 222210
rect 219206 212550 219266 222150
rect 219387 219332 219453 219333
rect 219387 219268 219388 219332
rect 219452 219268 219453 219332
rect 219387 219267 219453 219268
rect 219022 212490 219266 212550
rect 219022 122850 219082 212490
rect 219390 205650 219450 219267
rect 219206 205590 219450 205650
rect 219206 200130 219266 205590
rect 219206 200070 219450 200130
rect 219390 199610 219450 200070
rect 219206 199550 219450 199610
rect 219206 190770 219266 199550
rect 219206 190710 219450 190770
rect 219390 190470 219450 190710
rect 219206 190410 219450 190470
rect 219206 180810 219266 190410
rect 219206 180750 219450 180810
rect 219390 180570 219450 180750
rect 219206 180510 219450 180570
rect 219206 171730 219266 180510
rect 219206 171670 219634 171730
rect 219574 171150 219634 171670
rect 219206 171090 219634 171150
rect 219206 161490 219266 171090
rect 219206 161430 219634 161490
rect 219574 160850 219634 161430
rect 219206 160790 219634 160850
rect 219206 152010 219266 160790
rect 219206 151950 219450 152010
rect 219390 151830 219450 151950
rect 219206 151770 219450 151830
rect 219206 142170 219266 151770
rect 219206 142110 219450 142170
rect 219390 141810 219450 142110
rect 219206 141750 219450 141810
rect 219206 132970 219266 141750
rect 219206 132910 219450 132970
rect 219390 132510 219450 132910
rect 219206 132450 219450 132510
rect 219206 123450 219266 132450
rect 219206 123390 219634 123450
rect 219022 122790 219266 122850
rect 219019 121412 219085 121413
rect 219019 121348 219020 121412
rect 219084 121348 219085 121412
rect 219019 121347 219085 121348
rect 219022 118710 219082 121347
rect 219206 119645 219266 122790
rect 219574 121413 219634 123390
rect 219571 121412 219637 121413
rect 219571 121348 219572 121412
rect 219636 121348 219637 121412
rect 219571 121347 219637 121348
rect 219203 119644 219269 119645
rect 219203 119580 219204 119644
rect 219268 119580 219269 119644
rect 219203 119579 219269 119580
rect 219022 118650 219450 118710
rect 219390 113117 219450 118650
rect 219387 113116 219453 113117
rect 219387 113052 219388 113116
rect 219452 113052 219453 113116
rect 219387 113051 219453 113052
rect 220862 110941 220922 498067
rect 223619 337652 223685 337653
rect 223619 337588 223620 337652
rect 223684 337588 223685 337652
rect 223619 337587 223685 337588
rect 223622 118285 223682 337587
rect 224723 222460 224789 222461
rect 224723 222396 224724 222460
rect 224788 222396 224789 222460
rect 224723 222395 224789 222396
rect 224726 205650 224786 222395
rect 226931 220012 226997 220013
rect 226931 219948 226932 220012
rect 226996 219948 226997 220012
rect 226931 219947 226997 219948
rect 224726 205590 224970 205650
rect 224910 118710 224970 205590
rect 224910 118650 225154 118710
rect 223619 118284 223685 118285
rect 223619 118220 223620 118284
rect 223684 118220 223685 118284
rect 223619 118219 223685 118220
rect 223622 118013 223682 118219
rect 223619 118012 223685 118013
rect 223619 117948 223620 118012
rect 223684 117948 223685 118012
rect 223619 117947 223685 117948
rect 225094 112709 225154 118650
rect 226934 113117 226994 219947
rect 228590 119373 228650 606051
rect 230979 337380 231045 337381
rect 230979 337316 230980 337380
rect 231044 337316 231045 337380
rect 230979 337315 231045 337316
rect 228587 119372 228653 119373
rect 228587 119308 228588 119372
rect 228652 119308 228653 119372
rect 228587 119307 228653 119308
rect 228219 117468 228285 117469
rect 228219 117404 228220 117468
rect 228284 117404 228285 117468
rect 228219 117403 228285 117404
rect 226931 113116 226997 113117
rect 226931 113052 226932 113116
rect 226996 113052 226997 113116
rect 226931 113051 226997 113052
rect 225091 112708 225157 112709
rect 225091 112644 225092 112708
rect 225156 112644 225157 112708
rect 225091 112643 225157 112644
rect 220859 110940 220925 110941
rect 220859 110876 220860 110940
rect 220924 110876 220925 110940
rect 220859 110875 220925 110876
rect 222331 110532 222397 110533
rect 222331 110468 222332 110532
rect 222396 110468 222397 110532
rect 222331 110467 222397 110468
rect 222334 9213 222394 110467
rect 228222 10709 228282 117403
rect 228219 10708 228285 10709
rect 228219 10644 228220 10708
rect 228284 10644 228285 10708
rect 228219 10643 228285 10644
rect 230982 9213 231042 337315
rect 232454 111213 232514 616795
rect 233739 371788 233805 371789
rect 233739 371724 233740 371788
rect 233804 371724 233805 371788
rect 233739 371723 233805 371724
rect 232451 111212 232517 111213
rect 232451 111148 232452 111212
rect 232516 111148 232517 111212
rect 232451 111147 232517 111148
rect 233742 9485 233802 371723
rect 234662 118557 234722 616795
rect 243491 220012 243557 220013
rect 243491 219948 243492 220012
rect 243556 219948 243557 220012
rect 243491 219947 243557 219948
rect 240179 219740 240245 219741
rect 240179 219676 240180 219740
rect 240244 219676 240245 219740
rect 240179 219675 240245 219676
rect 235947 219468 236013 219469
rect 235947 219404 235948 219468
rect 236012 219404 236013 219468
rect 235947 219403 236013 219404
rect 234659 118556 234725 118557
rect 234659 118492 234660 118556
rect 234724 118492 234725 118556
rect 234659 118491 234725 118492
rect 235763 117468 235829 117469
rect 235763 117404 235764 117468
rect 235828 117404 235829 117468
rect 235763 117403 235829 117404
rect 235766 10709 235826 117403
rect 235950 111893 236010 219403
rect 240182 111893 240242 219675
rect 241651 117468 241717 117469
rect 241651 117404 241652 117468
rect 241716 117404 241717 117468
rect 241651 117403 241717 117404
rect 235947 111892 236013 111893
rect 235947 111828 235948 111892
rect 236012 111828 236013 111892
rect 235947 111827 236013 111828
rect 240179 111892 240245 111893
rect 240179 111828 240180 111892
rect 240244 111828 240245 111892
rect 240179 111827 240245 111828
rect 235763 10708 235829 10709
rect 235763 10644 235764 10708
rect 235828 10644 235829 10708
rect 235763 10643 235829 10644
rect 241654 10165 241714 117403
rect 241651 10164 241717 10165
rect 241651 10100 241652 10164
rect 241716 10100 241717 10164
rect 241651 10099 241717 10100
rect 233739 9484 233805 9485
rect 233739 9420 233740 9484
rect 233804 9420 233805 9484
rect 233739 9419 233805 9420
rect 222331 9212 222397 9213
rect 222331 9148 222332 9212
rect 222396 9148 222397 9212
rect 222331 9147 222397 9148
rect 230979 9212 231045 9213
rect 230979 9148 230980 9212
rect 231044 9148 231045 9212
rect 230979 9147 231045 9148
rect 212395 3772 212461 3773
rect 212395 3708 212396 3772
rect 212460 3708 212461 3772
rect 212395 3707 212461 3708
rect 217179 3772 217245 3773
rect 217179 3708 217180 3772
rect 217244 3708 217245 3772
rect 217179 3707 217245 3708
rect 190499 3636 190565 3637
rect 190499 3572 190500 3636
rect 190564 3572 190565 3636
rect 190499 3571 190565 3572
rect 243494 3501 243554 219947
rect 246254 118285 246314 616795
rect 258027 615636 258093 615637
rect 258027 615572 258028 615636
rect 258092 615572 258093 615636
rect 258027 615571 258093 615572
rect 258030 615510 258090 615571
rect 257846 615450 258090 615510
rect 248275 273868 248341 273869
rect 248275 273804 248276 273868
rect 248340 273804 248341 273868
rect 248275 273803 248341 273804
rect 246251 118284 246317 118285
rect 246251 118220 246252 118284
rect 246316 118220 246317 118284
rect 246251 118219 246317 118220
rect 248278 9485 248338 273803
rect 257846 224970 257906 615450
rect 283419 610060 283485 610061
rect 283419 609996 283420 610060
rect 283484 609996 283485 610060
rect 283419 609995 283485 609996
rect 268331 553484 268397 553485
rect 268331 553420 268332 553484
rect 268396 553420 268397 553484
rect 268331 553419 268397 553420
rect 276611 553484 276677 553485
rect 276611 553420 276612 553484
rect 276676 553420 276677 553484
rect 276611 553419 276677 553420
rect 263731 436116 263797 436117
rect 263731 436052 263732 436116
rect 263796 436052 263797 436116
rect 263731 436051 263797 436052
rect 263363 325004 263429 325005
rect 263363 324940 263364 325004
rect 263428 324940 263429 325004
rect 263363 324939 263429 324940
rect 261155 300932 261221 300933
rect 261155 300868 261156 300932
rect 261220 300868 261221 300932
rect 261155 300867 261221 300868
rect 257846 224910 258090 224970
rect 253059 220012 253125 220013
rect 253059 219948 253060 220012
rect 253124 219948 253125 220012
rect 253059 219947 253125 219948
rect 249011 118012 249077 118013
rect 249011 117948 249012 118012
rect 249076 117948 249077 118012
rect 249011 117947 249077 117948
rect 249014 10709 249074 117947
rect 253062 111893 253122 219947
rect 258030 215310 258090 224910
rect 257846 215250 258090 215310
rect 257846 128370 257906 215250
rect 261158 132510 261218 300867
rect 261158 132450 261402 132510
rect 257846 128310 258090 128370
rect 258030 120053 258090 128310
rect 258027 120052 258093 120053
rect 258027 119988 258028 120052
rect 258092 119988 258093 120052
rect 258027 119987 258093 119988
rect 261342 118693 261402 132450
rect 261339 118692 261405 118693
rect 261339 118628 261340 118692
rect 261404 118628 261405 118692
rect 261339 118627 261405 118628
rect 253979 118420 254045 118421
rect 253979 118356 253980 118420
rect 254044 118356 254045 118420
rect 253979 118355 254045 118356
rect 253059 111892 253125 111893
rect 253059 111828 253060 111892
rect 253124 111828 253125 111892
rect 253059 111827 253125 111828
rect 253982 10709 254042 118355
rect 261342 10709 261402 118627
rect 249011 10708 249077 10709
rect 249011 10644 249012 10708
rect 249076 10644 249077 10708
rect 249011 10643 249077 10644
rect 253979 10708 254045 10709
rect 253979 10644 253980 10708
rect 254044 10644 254045 10708
rect 253979 10643 254045 10644
rect 261339 10708 261405 10709
rect 261339 10644 261340 10708
rect 261404 10644 261405 10708
rect 261339 10643 261405 10644
rect 248275 9484 248341 9485
rect 248275 9420 248276 9484
rect 248340 9420 248341 9484
rect 248275 9419 248341 9420
rect 263366 4045 263426 324939
rect 263734 119373 263794 436051
rect 263731 119372 263797 119373
rect 263731 119308 263732 119372
rect 263796 119308 263797 119372
rect 263731 119307 263797 119308
rect 268334 9213 268394 553419
rect 274035 285700 274101 285701
rect 274035 285636 274036 285700
rect 274100 285636 274101 285700
rect 274035 285635 274101 285636
rect 273115 219468 273181 219469
rect 273115 219404 273116 219468
rect 273180 219404 273181 219468
rect 273115 219403 273181 219404
rect 269067 118148 269133 118149
rect 269067 118084 269068 118148
rect 269132 118084 269133 118148
rect 269067 118083 269133 118084
rect 269070 10709 269130 118083
rect 273118 113117 273178 219403
rect 273115 113116 273181 113117
rect 273115 113052 273116 113116
rect 273180 113052 273181 113116
rect 273115 113051 273181 113052
rect 274038 111077 274098 285635
rect 274035 111076 274101 111077
rect 274035 111012 274036 111076
rect 274100 111012 274101 111076
rect 274035 111011 274101 111012
rect 273667 110532 273733 110533
rect 273667 110468 273668 110532
rect 273732 110468 273733 110532
rect 273667 110467 273733 110468
rect 273670 10709 273730 110467
rect 269067 10708 269133 10709
rect 269067 10644 269068 10708
rect 269132 10644 269133 10708
rect 269067 10643 269133 10644
rect 273667 10708 273733 10709
rect 273667 10644 273668 10708
rect 273732 10644 273733 10708
rect 273667 10643 273733 10644
rect 276614 9621 276674 553419
rect 282683 432036 282749 432037
rect 282683 431972 282684 432036
rect 282748 431972 282749 432036
rect 282683 431971 282749 431972
rect 280659 220012 280725 220013
rect 280659 219948 280660 220012
rect 280724 219948 280725 220012
rect 280659 219947 280725 219948
rect 280662 111893 280722 219947
rect 282686 118965 282746 431971
rect 282683 118964 282749 118965
rect 282683 118900 282684 118964
rect 282748 118900 282749 118964
rect 282683 118899 282749 118900
rect 283422 117741 283482 609995
rect 289675 223684 289741 223685
rect 289675 223620 289676 223684
rect 289740 223620 289741 223684
rect 289675 223619 289741 223620
rect 283419 117740 283485 117741
rect 283419 117676 283420 117740
rect 283484 117676 283485 117740
rect 283419 117675 283485 117676
rect 282131 117468 282197 117469
rect 282131 117404 282132 117468
rect 282196 117404 282197 117468
rect 282131 117403 282197 117404
rect 280659 111892 280725 111893
rect 280659 111828 280660 111892
rect 280724 111828 280725 111892
rect 280659 111827 280725 111828
rect 282134 10709 282194 117403
rect 287099 117332 287165 117333
rect 287099 117268 287100 117332
rect 287164 117268 287165 117332
rect 287099 117267 287165 117268
rect 287102 10709 287162 117267
rect 282131 10708 282197 10709
rect 282131 10644 282132 10708
rect 282196 10644 282197 10708
rect 282131 10643 282197 10644
rect 287099 10708 287165 10709
rect 287099 10644 287100 10708
rect 287164 10644 287165 10708
rect 287099 10643 287165 10644
rect 276611 9620 276677 9621
rect 276611 9556 276612 9620
rect 276676 9556 276677 9620
rect 276611 9555 276677 9556
rect 268331 9212 268397 9213
rect 268331 9148 268332 9212
rect 268396 9148 268397 9212
rect 268331 9147 268397 9148
rect 289678 8533 289738 223619
rect 293171 219468 293237 219469
rect 293171 219404 293172 219468
rect 293236 219404 293237 219468
rect 293171 219403 293237 219404
rect 293174 111893 293234 219403
rect 295382 118557 295442 616795
rect 303291 249932 303357 249933
rect 303291 249868 303292 249932
rect 303356 249868 303357 249932
rect 303291 249867 303357 249868
rect 295379 118556 295445 118557
rect 295379 118492 295380 118556
rect 295444 118492 295445 118556
rect 295379 118491 295445 118492
rect 293907 117740 293973 117741
rect 293907 117676 293908 117740
rect 293972 117676 293973 117740
rect 293907 117675 293973 117676
rect 293171 111892 293237 111893
rect 293171 111828 293172 111892
rect 293236 111828 293237 111892
rect 293171 111827 293237 111828
rect 293910 109173 293970 117675
rect 303294 113933 303354 249867
rect 303291 113932 303357 113933
rect 303291 113868 303292 113932
rect 303356 113868 303357 113932
rect 303291 113867 303357 113868
rect 293907 109172 293973 109173
rect 293907 109108 293908 109172
rect 293972 109108 293973 109172
rect 293907 109107 293973 109108
rect 293910 10709 293970 109107
rect 293907 10708 293973 10709
rect 293907 10644 293908 10708
rect 293972 10644 293973 10708
rect 293907 10643 293973 10644
rect 289675 8532 289741 8533
rect 289675 8468 289676 8532
rect 289740 8468 289741 8532
rect 289675 8467 289741 8468
rect 263363 4044 263429 4045
rect 263363 3980 263364 4044
rect 263428 3980 263429 4044
rect 263363 3979 263429 3980
rect 243491 3500 243557 3501
rect 243491 3436 243492 3500
rect 243556 3436 243557 3500
rect 243491 3435 243557 3436
rect 138795 3228 138861 3229
rect 138795 3164 138796 3228
rect 138860 3164 138861 3228
rect 138795 3163 138861 3164
rect 119659 3092 119725 3093
rect 119659 3028 119660 3092
rect 119724 3028 119725 3092
rect 119659 3027 119725 3028
use sky130_fd_sc_hd__buf_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 35328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _352_
timestamp 1632766296
transform -1 0 65412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 78476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _397_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 78844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 77372 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 72036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _758_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 68816 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _462_
timestamp 1632766296
transform -1 0 88688 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _637_
timestamp 1632766296
transform 1 0 98624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _658_
timestamp 1632766296
transform 1 0 94944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 116932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _646_
timestamp 1632766296
transform -1 0 121440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _661_
timestamp 1632766296
transform 1 0 111504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _317_
timestamp 1632766296
transform -1 0 151432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _443_
timestamp 1632766296
transform 1 0 147660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _633_
timestamp 1632766296
transform -1 0 138276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _457_
timestamp 1632766296
transform -1 0 152812 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _734_
timestamp 1632766296
transform 1 0 168636 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _591_
timestamp 1632766296
transform -1 0 186024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _584_
timestamp 1632766296
transform 1 0 202860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471_
timestamp 1632766296
transform -1 0 225584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _272_
timestamp 1632766296
transform -1 0 244996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 248308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _468_
timestamp 1632766296
transform -1 0 240120 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1632766296
transform -1 0 277932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _604_
timestamp 1632766296
transform 1 0 261280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 270480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _745_
timestamp 1632766296
transform 1 0 272044 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _681_
timestamp 1632766296
transform -1 0 310868 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 335892 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _524_
timestamp 1632766296
transform 1 0 344448 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _356_
timestamp 1632766296
transform -1 0 456136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _687_
timestamp 1632766296
transform 1 0 478860 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1632766296
transform 1 0 496340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _301_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 9568 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _720_
timestamp 1632766296
transform 1 0 8004 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1632766296
transform 1 0 320344 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _588_
timestamp 1632766296
transform 1 0 310040 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _607_
timestamp 1632766296
transform 1 0 310040 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _690_
timestamp 1632766296
transform 1 0 310040 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_2  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 340584 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _586_
timestamp 1632766296
transform -1 0 346380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _777_
timestamp 1632766296
transform -1 0 343988 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _568_
timestamp 1632766296
transform -1 0 367080 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _609_
timestamp 1632766296
transform -1 0 376280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _728_
timestamp 1632766296
transform -1 0 373244 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _547_
timestamp 1632766296
transform 1 0 399280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _757_
timestamp 1632766296
transform -1 0 392380 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _579_
timestamp 1632766296
transform -1 0 408756 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _686_
timestamp 1632766296
transform 1 0 417864 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _762_
timestamp 1632766296
transform -1 0 416944 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _767_
timestamp 1632766296
transform -1 0 418968 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1632766296
transform 1 0 310040 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _578_
timestamp 1632766296
transform -1 0 310316 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _590_
timestamp 1632766296
transform -1 0 464140 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 3956 0 -1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _329_
timestamp 1632766296
transform 1 0 9292 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _354_
timestamp 1632766296
transform -1 0 9568 0 1 79424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _517_
timestamp 1632766296
transform 1 0 9292 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _595_
timestamp 1632766296
transform 1 0 7636 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _285_
timestamp 1632766296
transform -1 0 310316 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1632766296
transform -1 0 310316 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _454_
timestamp 1632766296
transform -1 0 338376 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 339388 0 1 78336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp 1632766296
transform -1 0 360364 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _288_
timestamp 1632766296
transform -1 0 372784 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _680_
timestamp 1632766296
transform 1 0 381708 0 -1 85952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _685_
timestamp 1632766296
transform 1 0 378396 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1632766296
transform -1 0 401304 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _556_
timestamp 1632766296
transform -1 0 394404 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _427_
timestamp 1632766296
transform 1 0 406088 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1632766296
transform 1 0 421912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _273_
timestamp 1632766296
transform 1 0 429640 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _733_
timestamp 1632766296
transform 1 0 438564 0 -1 90304
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _315_
timestamp 1632766296
transform 1 0 445372 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _420_
timestamp 1632766296
transform 1 0 442888 0 -1 79424
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _753_
timestamp 1632766296
transform -1 0 458252 0 1 99008
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _374_
timestamp 1632766296
transform 1 0 469292 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _516_
timestamp 1632766296
transform -1 0 477572 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _527_
timestamp 1632766296
transform 1 0 496248 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _531_
timestamp 1632766296
transform -1 0 494132 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _672_
timestamp 1632766296
transform -1 0 488152 0 -1 101184
box -38 -48 314 592
use SonarOnChip  soc1
timestamp 1633795376
transform 1 0 10000 0 1 10000
box 0 0 300000 100000
use sky130_fd_sc_hd__conb_1  _544_
timestamp 1632766296
transform 1 0 18768 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1632766296
transform -1 0 32660 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _437_
timestamp 1632766296
transform -1 0 35604 0 -1 119680
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _447_
timestamp 1632766296
transform 1 0 34500 0 1 118592
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _643_
timestamp 1632766296
transform 1 0 28244 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _673_
timestamp 1632766296
transform -1 0 33764 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1632766296
transform 1 0 38732 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _650_
timestamp 1632766296
transform -1 0 44068 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _656_
timestamp 1632766296
transform 1 0 50324 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _282_
timestamp 1632766296
transform -1 0 69460 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _419_
timestamp 1632766296
transform 1 0 63664 0 -1 119680
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _569_
timestamp 1632766296
transform 1 0 60996 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500_
timestamp 1632766296
transform 1 0 75348 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _526_
timestamp 1632766296
transform 1 0 81144 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _718_
timestamp 1632766296
transform 1 0 83076 0 -1 110976
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _494_
timestamp 1632766296
transform 1 0 102488 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _503_
timestamp 1632766296
transform -1 0 97152 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _611_
timestamp 1632766296
transform -1 0 101292 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _721_
timestamp 1632766296
transform 1 0 106444 0 -1 110976
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _542_
timestamp 1632766296
transform 1 0 131284 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _617_
timestamp 1632766296
transform 1 0 136988 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _466_
timestamp 1632766296
transform 1 0 145452 0 -1 119680
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1632766296
transform -1 0 170384 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _465_
timestamp 1632766296
transform -1 0 168452 0 -1 110976
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _554_
timestamp 1632766296
transform 1 0 172500 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _754_
timestamp 1632766296
transform -1 0 162472 0 -1 119680
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1632766296
transform 1 0 182620 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _446_
timestamp 1632766296
transform -1 0 179584 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _606_
timestamp 1632766296
transform 1 0 190256 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _743_
timestamp 1632766296
transform -1 0 180964 0 -1 110976
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_12  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 182988 0 1 110976
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 182252 0 -1 110976
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _277_
timestamp 1632766296
transform -1 0 209944 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _463_
timestamp 1632766296
transform 1 0 194304 0 -1 110976
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _549_
timestamp 1632766296
transform -1 0 202952 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _281_
timestamp 1632766296
transform 1 0 215464 0 -1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _359_
timestamp 1632766296
transform 1 0 221812 0 -1 110976
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _399_
timestamp 1632766296
transform -1 0 214728 0 -1 110976
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _513_
timestamp 1632766296
transform 1 0 224112 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _451_
timestamp 1632766296
transform 1 0 238464 0 -1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1632766296
transform -1 0 254380 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _648_
timestamp 1632766296
transform 1 0 248124 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _486_
timestamp 1632766296
transform 1 0 273424 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _679_
timestamp 1632766296
transform 1 0 273148 0 -1 110976
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _441_
timestamp 1632766296
transform -1 0 290628 0 -1 119680
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _535_
timestamp 1632766296
transform 1 0 286028 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492_
timestamp 1632766296
transform 1 0 307832 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _707_
timestamp 1632766296
transform -1 0 327796 0 -1 112064
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer16
timestamp 1632766296
transform -1 0 328808 0 1 110976
box -38 -48 682 592
use sky130_fd_sc_hd__buf_12  rebuffer17
timestamp 1632766296
transform -1 0 329636 0 -1 112064
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  rebuffer18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 328716 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _448_
timestamp 1632766296
transform -1 0 368644 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _284_
timestamp 1632766296
transform 1 0 419336 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _406_
timestamp 1632766296
transform -1 0 453284 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _581_
timestamp 1632766296
transform -1 0 440588 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _781_
timestamp 1632766296
transform -1 0 451720 0 -1 117504
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _533_
timestamp 1632766296
transform -1 0 457240 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _566_
timestamp 1632766296
transform -1 0 485484 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _567_
timestamp 1632766296
transform 1 0 480424 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518_
timestamp 1632766296
transform -1 0 496616 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1632766296
transform 1 0 9292 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _353_
timestamp 1632766296
transform 1 0 4508 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _407_
timestamp 1632766296
transform -1 0 9568 0 1 132736
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _483_
timestamp 1632766296
transform 1 0 7084 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _583_
timestamp 1632766296
transform 1 0 310040 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _380_
timestamp 1632766296
transform -1 0 367448 0 1 122944
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _540_
timestamp 1632766296
transform 1 0 356500 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _634_
timestamp 1632766296
transform 1 0 355764 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _655_
timestamp 1632766296
transform -1 0 383916 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _299_
timestamp 1632766296
transform -1 0 429640 0 -1 125120
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1632766296
transform 1 0 477664 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475_
timestamp 1632766296
transform 1 0 9292 0 -1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _309_
timestamp 1632766296
transform 1 0 321356 0 -1 152320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _662_
timestamp 1632766296
transform -1 0 315744 0 -1 147968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 321448 0 1 152320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer29
timestamp 1632766296
transform -1 0 323656 0 1 152320
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  _640_
timestamp 1632766296
transform 1 0 357144 0 1 147968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _537_
timestamp 1632766296
transform -1 0 389620 0 -1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _752_
timestamp 1632766296
transform 1 0 416116 0 1 140352
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _670_
timestamp 1632766296
transform -1 0 427524 0 -1 152320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _577_
timestamp 1632766296
transform -1 0 457976 0 -1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _644_
timestamp 1632766296
transform -1 0 455216 0 1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _268_
timestamp 1632766296
transform 1 0 9292 0 1 203456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1632766296
transform -1 0 8280 0 1 156672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _774_
timestamp 1632766296
transform -1 0 5060 0 1 169728
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _278_
timestamp 1632766296
transform 1 0 310040 0 -1 178432
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp 1632766296
transform 1 0 310040 0 -1 176256
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 310040 0 -1 202368
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _416_
timestamp 1632766296
transform -1 0 310776 0 -1 183872
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _715_
timestamp 1632766296
transform -1 0 336628 0 -1 176256
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer15
timestamp 1632766296
transform 1 0 336996 0 -1 176256
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 385848 0 -1 162112
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  _623_
timestamp 1632766296
transform -1 0 397716 0 1 194752
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _678_
timestamp 1632766296
transform 1 0 380696 0 -1 162112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _271_
timestamp 1632766296
transform -1 0 407652 0 1 179520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _558_
timestamp 1632766296
transform -1 0 415104 0 -1 162112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _632_
timestamp 1632766296
transform -1 0 414000 0 -1 201280
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer31
timestamp 1632766296
transform 1 0 406364 0 1 179520
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _487_
timestamp 1632766296
transform -1 0 466256 0 -1 162112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _585_
timestamp 1632766296
transform -1 0 450800 0 -1 195840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _504_
timestamp 1632766296
transform -1 0 484104 0 -1 200192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _541_
timestamp 1632766296
transform 1 0 484012 0 1 156672
box -38 -48 314 592
use SonarOnChip  soc2
timestamp 1633795376
transform 1 0 10000 0 1 120000
box 0 0 300000 100000
use sky130_fd_sc_hd__conb_1  _598_
timestamp 1632766296
transform 1 0 3036 0 -1 209984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _660_
timestamp 1632766296
transform 1 0 54832 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1632766296
transform -1 0 50140 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _682_
timestamp 1632766296
transform -1 0 79856 0 -1 220864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _667_
timestamp 1632766296
transform 1 0 77556 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1632766296
transform -1 0 75808 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _694_
timestamp 1632766296
transform -1 0 97152 0 -1 220864
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1632766296
transform -1 0 101016 0 1 224128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _740_
timestamp 1632766296
transform -1 0 133308 0 -1 220864
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _701_
timestamp 1632766296
transform -1 0 130088 0 -1 220864
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1632766296
transform -1 0 123556 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _741_
timestamp 1632766296
transform 1 0 162748 0 -1 220864
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1632766296
transform 1 0 178296 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _355_
timestamp 1632766296
transform 1 0 204976 0 -1 220864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _564_
timestamp 1632766296
transform 1 0 227700 0 1 223040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _555_
timestamp 1632766296
transform 1 0 235060 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _772_
timestamp 1632766296
transform -1 0 266524 0 -1 220864
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _371_
timestamp 1632766296
transform -1 0 257876 0 -1 220864
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 259624 0 -1 220864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _292_
timestamp 1632766296
transform 1 0 260452 0 1 223040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _575_
timestamp 1632766296
transform -1 0 288512 0 -1 220864
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer14
timestamp 1632766296
transform -1 0 290352 0 -1 225216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _698_
timestamp 1632766296
transform -1 0 290076 0 1 224128
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _654_
timestamp 1632766296
transform -1 0 310316 0 1 209984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _576_
timestamp 1632766296
transform 1 0 346840 0 1 225216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _485_
timestamp 1632766296
transform -1 0 346104 0 -1 218688
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _296_
timestamp 1632766296
transform -1 0 371864 0 1 216512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp 1632766296
transform 1 0 20332 0 1 237184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _778_
timestamp 1632766296
transform 1 0 61088 0 1 236096
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _565_
timestamp 1632766296
transform 1 0 115000 0 -1 244800
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4
timestamp 1632766296
transform -1 0 137264 0 -1 227392
box -38 -48 682 592
use sky130_fd_sc_hd__buf_12  rebuffer3
timestamp 1632766296
transform 1 0 136252 0 1 227392
box -38 -48 1510 592
use sky130_fd_sc_hd__o221a_2  _426_
timestamp 1632766296
transform -1 0 136252 0 -1 227392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1632766296
transform 1 0 153364 0 1 229568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _703_
timestamp 1632766296
transform -1 0 167900 0 -1 228480
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636_
timestamp 1632766296
transform 1 0 216016 0 -1 231744
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _573_
timestamp 1632766296
transform -1 0 240580 0 -1 232832
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _631_
timestamp 1632766296
transform 1 0 292008 0 -1 228480
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _523_
timestamp 1632766296
transform 1 0 315560 0 1 240448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _770_
timestamp 1632766296
transform -1 0 342608 0 1 236096
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _677_
timestamp 1632766296
transform 1 0 418508 0 1 230656
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _348_
timestamp 1632766296
transform 1 0 430744 0 1 237184
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 467360 0 1 240448
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _630_
timestamp 1632766296
transform 1 0 36156 0 -1 266560
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _559_
timestamp 1632766296
transform 1 0 59800 0 1 258944
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _747_
timestamp 1632766296
transform 1 0 77832 0 -1 264384
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _615_
timestamp 1632766296
transform 1 0 98532 0 -1 264384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _287_
timestamp 1632766296
transform -1 0 92552 0 1 269824
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _385_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 125304 0 -1 261120
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _293_
timestamp 1632766296
transform -1 0 118036 0 1 252416
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _580_
timestamp 1632766296
transform -1 0 139288 0 1 252416
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _683_
timestamp 1632766296
transform -1 0 181332 0 1 258944
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _732_
timestamp 1632766296
transform -1 0 220616 0 1 254592
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _460_
timestamp 1632766296
transform 1 0 207092 0 1 262208
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _739_
timestamp 1632766296
transform 1 0 230920 0 -1 251328
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _280_
timestamp 1632766296
transform 1 0 228712 0 1 267648
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _440_
timestamp 1632766296
transform -1 0 303232 0 -1 250240
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _294_
timestamp 1632766296
transform -1 0 299552 0 -1 256768
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _594_
timestamp 1632766296
transform 1 0 314916 0 -1 249152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1632766296
transform -1 0 317860 0 1 260032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _497_
timestamp 1632766296
transform -1 0 353648 0 1 265472
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _303_
timestamp 1632766296
transform -1 0 367540 0 1 266560
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _665_
timestamp 1632766296
transform 1 0 396428 0 1 254592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _639_
timestamp 1632766296
transform -1 0 380880 0 -1 254592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _657_
timestamp 1632766296
transform -1 0 442520 0 1 265472
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _714_
timestamp 1632766296
transform 1 0 443624 0 -1 252416
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _773_
timestamp 1632766296
transform -1 0 487048 0 1 266560
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1632766296
transform 1 0 470488 0 1 256768
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _308_
timestamp 1632766296
transform 1 0 483552 0 -1 257856
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _551_
timestamp 1632766296
transform 1 0 16652 0 1 281792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490_
timestamp 1632766296
transform -1 0 84824 0 -1 281792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _318_
timestamp 1632766296
transform -1 0 93196 0 -1 288320
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _729_
timestamp 1632766296
transform 1 0 137908 0 -1 292672
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _664_
timestamp 1632766296
transform 1 0 176732 0 1 277440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _386_
timestamp 1632766296
transform 1 0 158700 0 -1 274176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _750_
timestamp 1632766296
transform 1 0 243064 0 -1 283968
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _589_
timestamp 1632766296
transform -1 0 229356 0 1 273088
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _761_
timestamp 1632766296
transform 1 0 264316 0 -1 279616
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1632766296
transform -1 0 248768 0 -1 276352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _398_
timestamp 1632766296
transform 1 0 273608 0 -1 287232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  rebuffer7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 296332 0 1 282880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 297620 0 -1 283968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  rebuffer5
timestamp 1632766296
transform 1 0 296700 0 1 282880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  rebuffer10
timestamp 1632766296
transform 1 0 296700 0 -1 282880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _300_
timestamp 1632766296
transform 1 0 296056 0 -1 282880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1632766296
transform -1 0 329820 0 -1 280704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _360_
timestamp 1632766296
transform -1 0 341504 0 -1 291584
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer33
timestamp 1632766296
transform -1 0 374348 0 -1 270912
box -38 -48 682 592
use sky130_fd_sc_hd__buf_12  rebuffer30
timestamp 1632766296
transform 1 0 373704 0 1 270912
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _270_
timestamp 1632766296
transform 1 0 373060 0 1 270912
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _501_
timestamp 1632766296
transform -1 0 420808 0 -1 273088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _612_
timestamp 1632766296
transform 1 0 482816 0 1 282880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _766_
timestamp 1632766296
transform -1 0 6164 0 -1 304640
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _563_
timestamp 1632766296
transform -1 0 46736 0 1 298112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477_
timestamp 1632766296
transform 1 0 83996 0 1 292672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481_
timestamp 1632766296
transform 1 0 104328 0 1 293760
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _351_
timestamp 1632766296
transform 1 0 111964 0 -1 295936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _748_
timestamp 1632766296
transform -1 0 262568 0 1 301376
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _562_
timestamp 1632766296
transform 1 0 274528 0 -1 293760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _519_
timestamp 1632766296
transform -1 0 326048 0 -1 303552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _306_
timestamp 1632766296
transform 1 0 340860 0 -1 301376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _393_
timestamp 1632766296
transform 1 0 414184 0 1 295936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _713_
timestamp 1632766296
transform -1 0 22172 0 1 305728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _676_
timestamp 1632766296
transform -1 0 21528 0 -1 317696
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _744_
timestamp 1632766296
transform 1 0 50048 0 1 304640
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _572_
timestamp 1632766296
transform 1 0 78752 0 -1 319872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478_
timestamp 1632766296
transform 1 0 91356 0 -1 326400
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _297_
timestamp 1632766296
transform 1 0 93288 0 -1 326400
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _695_
timestamp 1632766296
transform -1 0 141312 0 1 306816
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _724_
timestamp 1632766296
transform -1 0 184828 0 -1 312256
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _512_
timestamp 1632766296
transform 1 0 187220 0 -1 306816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _495_
timestamp 1632766296
transform 1 0 181884 0 -1 317696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _560_
timestamp 1632766296
transform -1 0 282532 0 -1 325312
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _722_
timestamp 1632766296
transform -1 0 342332 0 1 318784
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _626_
timestamp 1632766296
transform 1 0 348220 0 -1 323136
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _401_
timestamp 1632766296
transform 1 0 331568 0 -1 325312
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _529_
timestamp 1632766296
transform -1 0 403604 0 -1 311168
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _324_
timestamp 1632766296
transform -1 0 427248 0 -1 308992
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _506_
timestamp 1632766296
transform -1 0 450800 0 1 325312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _548_
timestamp 1632766296
transform -1 0 465704 0 1 319872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1632766296
transform 1 0 481712 0 -1 314432
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _332_
timestamp 1632766296
transform -1 0 9936 0 1 332928
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _613_
timestamp 1632766296
transform 1 0 29348 0 1 343808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _649_
timestamp 1632766296
transform 1 0 62008 0 -1 332928
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _491_
timestamp 1632766296
transform 1 0 67988 0 1 335104
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _601_
timestamp 1632766296
transform -1 0 87308 0 1 326400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472_
timestamp 1632766296
transform 1 0 87584 0 -1 331840
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _768_
timestamp 1632766296
transform -1 0 106444 0 -1 336192
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _502_
timestamp 1632766296
transform -1 0 208748 0 1 327488
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 219052 0 1 337280
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _696_
timestamp 1632766296
transform -1 0 233404 0 1 343808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _493_
timestamp 1632766296
transform -1 0 252632 0 -1 329664
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _381_
timestamp 1632766296
transform -1 0 311236 0 1 334016
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _314_
timestamp 1632766296
transform 1 0 344540 0 -1 339456
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _610_
timestamp 1632766296
transform -1 0 366068 0 -1 335104
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _561_
timestamp 1632766296
transform 1 0 363308 0 1 330752
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479_
timestamp 1632766296
transform -1 0 376464 0 -1 344896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _433_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 381248 0 -1 329664
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1632766296
transform 1 0 385112 0 -1 338368
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _608_
timestamp 1632766296
transform -1 0 411240 0 1 339456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1632766296
transform 1 0 423936 0 -1 327488
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 438288 0 -1 329664
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _339_
timestamp 1632766296
transform 1 0 485392 0 -1 347072
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _418_
timestamp 1632766296
transform -1 0 5336 0 1 348160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1632766296
transform -1 0 7544 0 1 355776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _499_
timestamp 1632766296
transform 1 0 49680 0 1 362304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _775_
timestamp 1632766296
transform 1 0 89240 0 -1 356864
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _295_
timestamp 1632766296
transform -1 0 88412 0 1 359040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _625_
timestamp 1632766296
transform 1 0 140852 0 1 351424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _430_
timestamp 1632766296
transform -1 0 143428 0 -1 365568
box -38 -48 498 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 1632766296
transform -1 0 194212 0 1 353600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_12  rebuffer8
timestamp 1632766296
transform -1 0 196052 0 1 353600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  rebuffer28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 195500 0 -1 353600
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer27
timestamp 1632766296
transform -1 0 195132 0 -1 354688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _307_
timestamp 1632766296
transform 1 0 193292 0 -1 353600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _261_
timestamp 1632766296
transform -1 0 180504 0 1 362304
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _629_
timestamp 1632766296
transform -1 0 200284 0 1 355776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _635_
timestamp 1632766296
transform 1 0 244168 0 1 360128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1632766296
transform 1 0 293664 0 1 368832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _435_
timestamp 1632766296
transform -1 0 361652 0 1 355776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _346_
timestamp 1632766296
transform 1 0 361468 0 -1 360128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _310_
timestamp 1632766296
transform 1 0 360180 0 -1 366656
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _616_
timestamp 1632766296
transform -1 0 403972 0 -1 355776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _458_
timestamp 1632766296
transform 1 0 402776 0 1 360128
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1632766296
transform 1 0 451444 0 1 349248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _782_
timestamp 1632766296
transform 1 0 470396 0 1 364480
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1632766296
transform 1 0 473616 0 -1 365568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _736_
timestamp 1632766296
transform -1 0 40848 0 1 380800
box -38 -48 1602 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer22
timestamp 1632766296
transform -1 0 72036 0 1 378624
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _442_
timestamp 1632766296
transform -1 0 70932 0 1 378624
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_2  _392_
timestamp 1632766296
transform 1 0 88780 0 1 384064
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _620_
timestamp 1632766296
transform -1 0 96600 0 1 382976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _602_
timestamp 1632766296
transform 1 0 108100 0 -1 385152
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _467_
timestamp 1632766296
transform 1 0 103224 0 1 384064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _275_
timestamp 1632766296
transform -1 0 96048 0 1 374272
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _521_
timestamp 1632766296
transform -1 0 130640 0 1 382976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _349_
timestamp 1632766296
transform -1 0 132664 0 1 384064
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _286_
timestamp 1632766296
transform 1 0 176916 0 -1 384064
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _702_
timestamp 1632766296
transform 1 0 199548 0 -1 384064
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _675_
timestamp 1632766296
transform 1 0 214544 0 1 369920
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _508_
timestamp 1632766296
transform -1 0 207828 0 1 375360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1632766296
transform 1 0 233680 0 -1 372096
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _659_
timestamp 1632766296
transform -1 0 274712 0 -1 380800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _756_
timestamp 1632766296
transform 1 0 308292 0 1 375360
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _628_
timestamp 1632766296
transform -1 0 322552 0 1 382976
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _283_
timestamp 1632766296
transform 1 0 346196 0 1 387328
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _453_
timestamp 1632766296
transform -1 0 368184 0 -1 387328
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _717_
timestamp 1632766296
transform 1 0 409032 0 -1 375360
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _511_
timestamp 1632766296
transform -1 0 442244 0 1 372096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _274_
timestamp 1632766296
transform -1 0 450708 0 1 374272
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476_
timestamp 1632766296
transform -1 0 20792 0 -1 393856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _429_
timestamp 1632766296
transform 1 0 11776 0 1 394944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _305_
timestamp 1632766296
transform -1 0 23092 0 -1 394944
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _520_
timestamp 1632766296
transform 1 0 42872 0 -1 396032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _553_
timestamp 1632766296
transform -1 0 56856 0 -1 403648
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _365_
timestamp 1632766296
transform -1 0 67804 0 1 400384
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _505_
timestamp 1632766296
transform -1 0 170200 0 1 401472
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484_
timestamp 1632766296
transform 1 0 256864 0 -1 392768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp 1632766296
transform 1 0 252908 0 1 399296
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _627_
timestamp 1632766296
transform 1 0 282440 0 1 396032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _545_
timestamp 1632766296
transform 1 0 268732 0 -1 400384
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _603_
timestamp 1632766296
transform -1 0 313996 0 -1 396032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509_
timestamp 1632766296
transform -1 0 326784 0 -1 398208
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _552_
timestamp 1632766296
transform -1 0 341044 0 1 397120
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _322_
timestamp 1632766296
transform 1 0 380512 0 1 394944
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _536_
timestamp 1632766296
transform 1 0 399832 0 1 398208
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _704_
timestamp 1632766296
transform 1 0 451536 0 1 393856
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _414_
timestamp 1632766296
transform 1 0 27416 0 -1 423232
box -38 -48 958 592
use sky130_fd_sc_hd__or2_2  _404_
timestamp 1632766296
transform -1 0 55752 0 -1 410176
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _289_
timestamp 1632766296
transform 1 0 56580 0 1 409088
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _622_
timestamp 1632766296
transform 1 0 113896 0 -1 405824
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _600_
timestamp 1632766296
transform 1 0 119416 0 1 414528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _445_
timestamp 1632766296
transform 1 0 112424 0 1 410176
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _394_
timestamp 1632766296
transform 1 0 99636 0 -1 411264
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _618_
timestamp 1632766296
transform 1 0 136344 0 1 416704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _596_
timestamp 1632766296
transform 1 0 143612 0 1 412352
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _361_
timestamp 1632766296
transform 1 0 133676 0 1 423232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _474_
timestamp 1632766296
transform 1 0 151248 0 -1 412352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 1632766296
transform -1 0 239384 0 1 424320
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _755_
timestamp 1632766296
transform -1 0 260360 0 1 413440
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _699_
timestamp 1632766296
transform 1 0 256496 0 -1 415616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _276_
timestamp 1632766296
transform 1 0 278944 0 -1 415616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _668_
timestamp 1632766296
transform -1 0 338652 0 1 411264
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _391_
timestamp 1632766296
transform 1 0 331108 0 1 423232
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _291_
timestamp 1632766296
transform 1 0 333684 0 -1 417792
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _759_
timestamp 1632766296
transform 1 0 402408 0 -1 414528
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _449_
timestamp 1632766296
transform -1 0 412712 0 -1 428672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _719_
timestamp 1632766296
transform -1 0 443992 0 1 421056
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _488_
timestamp 1632766296
transform -1 0 442060 0 1 405824
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482_
timestamp 1632766296
transform -1 0 450800 0 1 426496
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer26
timestamp 1632766296
transform 1 0 42412 0 -1 439552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  rebuffer25
timestamp 1632766296
transform 1 0 42412 0 1 439552
box -38 -48 1510 592
use sky130_fd_sc_hd__o311a_2  _434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform 1 0 47472 0 -1 435200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _298_
timestamp 1632766296
transform 1 0 41768 0 -1 439552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _653_
timestamp 1632766296
transform 1 0 64584 0 -1 448256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514_
timestamp 1632766296
transform 1 0 63848 0 1 433024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489_
timestamp 1632766296
transform -1 0 57040 0 -1 435200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _304_
timestamp 1632766296
transform 1 0 53360 0 -1 451520
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _396_
timestamp 1632766296
transform -1 0 91908 0 1 434112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _705_
timestamp 1632766296
transform 1 0 111872 0 -1 447168
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _330_
timestamp 1632766296
transform 1 0 142232 0 -1 429760
box -38 -48 498 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer21
timestamp 1632766296
transform 1 0 152352 0 1 442816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer20
timestamp 1632766296
transform -1 0 153916 0 -1 443904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _700_
timestamp 1632766296
transform 1 0 151984 0 -1 443904
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_2  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1632766296
transform -1 0 176364 0 1 448256
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _725_
timestamp 1632766296
transform 1 0 281336 0 1 431936
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _587_
timestamp 1632766296
transform 1 0 281152 0 -1 442816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _769_
timestamp 1632766296
transform -1 0 334972 0 -1 447168
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1632766296
transform -1 0 376280 0 1 441728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _557_
timestamp 1632766296
transform -1 0 397348 0 -1 437376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _452_
timestamp 1632766296
transform -1 0 419152 0 1 439552
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1632766296
transform 1 0 423936 0 -1 443904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _710_
timestamp 1632766296
transform 1 0 93380 0 1 473280
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _570_
timestamp 1632766296
transform -1 0 110032 0 -1 463488
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _444_
timestamp 1632766296
transform 1 0 111780 0 1 466752
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _528_
timestamp 1632766296
transform 1 0 133584 0 -1 454784
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _735_
timestamp 1632766296
transform 1 0 149316 0 -1 471104
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _543_
timestamp 1632766296
transform 1 0 170200 0 -1 461312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _532_
timestamp 1632766296
transform 1 0 185380 0 -1 458048
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _751_
timestamp 1632766296
transform 1 0 194764 0 1 466752
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_2  _431_
timestamp 1632766296
transform -1 0 198720 0 1 471104
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _290_
timestamp 1632766296
transform 1 0 202676 0 1 473280
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  rebuffer19
timestamp 1632766296
transform -1 0 224572 0 -1 465664
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _691_
timestamp 1632766296
transform 1 0 222640 0 -1 465664
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1632766296
transform -1 0 254288 0 1 456960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538_
timestamp 1632766296
transform -1 0 315560 0 -1 453696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _571_
timestamp 1632766296
transform -1 0 363032 0 1 463488
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _737_
timestamp 1632766296
transform 1 0 432492 0 -1 470016
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_2  _312_
timestamp 1632766296
transform -1 0 495972 0 1 475456
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _712_
timestamp 1632766296
transform -1 0 21528 0 -1 487424
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _316_
timestamp 1632766296
transform -1 0 16652 0 -1 480896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _697_
timestamp 1632766296
transform -1 0 32844 0 1 492864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _621_
timestamp 1632766296
transform -1 0 190624 0 -1 500480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _771_
timestamp 1632766296
transform -1 0 208564 0 1 491776
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _666_
timestamp 1632766296
transform -1 0 205160 0 -1 495040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _400_
timestamp 1632766296
transform -1 0 208656 0 -1 498304
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _749_
timestamp 1632766296
transform 1 0 238188 0 1 479808
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _496_
timestamp 1632766296
transform -1 0 229356 0 1 493952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  rebuffer23
timestamp 1632766296
transform 1 0 255576 0 1 496128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  rebuffer13
timestamp 1632766296
transform 1 0 256312 0 -1 496128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  rebuffer12
timestamp 1632766296
transform 1 0 256312 0 1 496128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _779_
timestamp 1632766296
transform 1 0 248032 0 1 489600
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_2  _341_
timestamp 1632766296
transform -1 0 264132 0 1 485248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp 1632766296
transform 1 0 255668 0 -1 496128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _746_
timestamp 1632766296
transform 1 0 276920 0 1 491776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _764_
timestamp 1632766296
transform -1 0 384008 0 1 481984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _742_
timestamp 1632766296
transform 1 0 412896 0 1 489600
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _439_
timestamp 1632766296
transform -1 0 418232 0 -1 487424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _546_
timestamp 1632766296
transform -1 0 470304 0 -1 489600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _423_
timestamp 1632766296
transform -1 0 464600 0 -1 484160
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _642_
timestamp 1632766296
transform 1 0 116564 0 -1 502656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1632766296
transform -1 0 384008 0 -1 504832
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_2  _342_
timestamp 1632766296
transform -1 0 421360 0 1 500480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _730_
timestamp 1632766296
transform -1 0 13064 0 1 527680
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _614_
timestamp 1632766296
transform 1 0 24196 0 1 513536
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _411_
timestamp 1632766296
transform -1 0 11776 0 1 524416
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _258_
timestamp 1632766296
transform -1 0 46276 0 1 513536
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _480_
timestamp 1632766296
transform -1 0 91632 0 -1 528768
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1632766296
transform 1 0 92000 0 -1 514624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1632766296
transform -1 0 121164 0 -1 526592
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer35
timestamp 1632766296
transform -1 0 249320 0 -1 507008
box -38 -48 682 592
use sky130_fd_sc_hd__buf_12  rebuffer34
timestamp 1632766296
transform -1 0 250148 0 1 507008
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_2  _470_
timestamp 1632766296
transform -1 0 248308 0 1 507008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _776_
timestamp 1632766296
transform -1 0 260728 0 1 513536
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _692_
timestamp 1632766296
transform -1 0 263212 0 -1 525504
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _716_
timestamp 1632766296
transform 1 0 290720 0 -1 518976
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _763_
timestamp 1632766296
transform 1 0 324944 0 -1 508096
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _624_
timestamp 1632766296
transform 1 0 317124 0 -1 511360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1632766296
transform -1 0 319976 0 1 514624
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer24
timestamp 1632766296
transform 1 0 351440 0 -1 525504
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _693_
timestamp 1632766296
transform 1 0 351072 0 1 524416
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _525_
timestamp 1632766296
transform 1 0 353740 0 1 527680
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1632766296
transform -1 0 355672 0 1 528768
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _726_
timestamp 1632766296
transform -1 0 377108 0 -1 527680
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _708_
timestamp 1632766296
transform 1 0 405352 0 -1 514624
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _262_
timestamp 1632766296
transform 1 0 426604 0 -1 508096
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _515_
timestamp 1632766296
transform -1 0 17572 0 1 537472
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _319_
timestamp 1632766296
transform 1 0 59064 0 -1 539648
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _473_
timestamp 1632766296
transform 1 0 121624 0 -1 547264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _450_
timestamp 1632766296
transform 1 0 119416 0 -1 541824
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1632766296
transform -1 0 136252 0 -1 534208
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _464_
timestamp 1632766296
transform 1 0 157228 0 -1 544000
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _413_
timestamp 1632766296
transform 1 0 158424 0 -1 540736
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _780_
timestamp 1632766296
transform 1 0 231840 0 1 548352
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_2  _267_
timestamp 1632766296
transform -1 0 268916 0 -1 553792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _669_
timestamp 1632766296
transform 1 0 304704 0 1 554880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _597_
timestamp 1632766296
transform -1 0 328164 0 1 536384
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _539_
timestamp 1632766296
transform 1 0 330648 0 1 553792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _455_
timestamp 1632766296
transform 1 0 331292 0 1 534208
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522_
timestamp 1632766296
transform -1 0 342700 0 -1 532032
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _723_
timestamp 1632766296
transform -1 0 380696 0 1 547264
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _651_
timestamp 1632766296
transform -1 0 416852 0 1 544000
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _357_
timestamp 1632766296
transform -1 0 435436 0 1 551616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _663_
timestamp 1632766296
transform -1 0 442152 0 1 537472
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _605_
timestamp 1632766296
transform -1 0 445280 0 1 544000
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _390_
timestamp 1632766296
transform 1 0 14904 0 1 561408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _592_
timestamp 1632766296
transform 1 0 78384 0 1 565760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _410_
timestamp 1632766296
transform 1 0 75624 0 1 565760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _574_
timestamp 1632766296
transform 1 0 113436 0 1 578816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _456_
timestamp 1632766296
transform -1 0 170200 0 -1 557056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _765_
timestamp 1632766296
transform 1 0 196420 0 -1 572288
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _320_
timestamp 1632766296
transform -1 0 204424 0 -1 559232
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _731_
timestamp 1632766296
transform -1 0 237912 0 -1 571200
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _599_
timestamp 1632766296
transform -1 0 248492 0 -1 578816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _671_
timestamp 1632766296
transform 1 0 285108 0 -1 571200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _395_
timestamp 1632766296
transform -1 0 325956 0 1 565760
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _619_
timestamp 1632766296
transform -1 0 369656 0 -1 572288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507_
timestamp 1632766296
transform -1 0 376740 0 1 569024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _706_
timestamp 1632766296
transform 1 0 402868 0 1 557056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _689_
timestamp 1632766296
transform 1 0 396244 0 1 578816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _550_
timestamp 1632766296
transform -1 0 417772 0 -1 576640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _469_
timestamp 1632766296
transform 1 0 423384 0 1 576640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _711_
timestamp 1632766296
transform 1 0 482172 0 -1 580992
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _459_
timestamp 1632766296
transform 1 0 473708 0 1 566848
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _760_
timestamp 1632766296
transform 1 0 22724 0 1 600576
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _368_
timestamp 1632766296
transform -1 0 50784 0 -1 599488
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _534_
timestamp 1632766296
transform 1 0 106536 0 1 584256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _688_
timestamp 1632766296
transform 1 0 205436 0 1 596224
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _684_
timestamp 1632766296
transform -1 0 202032 0 -1 584256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _647_
timestamp 1632766296
transform 1 0 184368 0 -1 601664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _638_
timestamp 1632766296
transform 1 0 233220 0 -1 600576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _582_
timestamp 1632766296
transform 1 0 247388 0 1 596224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _645_
timestamp 1632766296
transform -1 0 322460 0 1 603840
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _641_
timestamp 1632766296
transform 1 0 313168 0 -1 586432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _652_
timestamp 1632766296
transform 1 0 405720 0 1 583168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498_
timestamp 1632766296
transform -1 0 410596 0 1 585344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _421_
timestamp 1632766296
transform 1 0 419336 0 -1 590784
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _321_
timestamp 1632766296
transform -1 0 463864 0 -1 587520
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _727_
timestamp 1632766296
transform -1 0 494408 0 1 590784
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1632766296
transform -1 0 200560 0 1 607104
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _358_
timestamp 1632766296
transform 1 0 282992 0 1 610368
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _424_
timestamp 1632766296
transform -1 0 168084 0 1 613632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _438_
timestamp 1632766296
transform -1 0 376280 0 1 611456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _461_
timestamp 1632766296
transform -1 0 334972 0 -1 608192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _510_
timestamp 1632766296
transform 1 0 129444 0 -1 609280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _593_
timestamp 1632766296
transform 1 0 200652 0 1 609280
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _674_
timestamp 1632766296
transform 1 0 364044 0 1 614720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _738_
timestamp 1632766296
transform 1 0 228160 0 -1 607104
box -38 -48 1602 592
<< labels >>
rlabel metal2 s 451158 -960 451270 480 8 io_in[0]
port 0 nsew signal input
rlabel metal2 s 27222 -960 27334 480 8 io_in[10]
port 1 nsew signal input
rlabel metal3 s 499520 245836 500960 246076 6 io_in[11]
port 2 nsew signal input
rlabel metal3 s -960 147644 480 147884 4 io_in[12]
port 3 nsew signal input
rlabel metal2 s 189326 619520 189438 620960 6 io_in[13]
port 4 nsew signal input
rlabel metal3 s 499520 389180 500960 389420 6 io_in[14]
port 5 nsew signal input
rlabel metal2 s 165222 619520 165334 620960 6 io_in[15]
port 6 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[16]
port 7 nsew signal input
rlabel metal3 s 499520 590732 500960 590972 6 io_in[17]
port 8 nsew signal input
rlabel metal3 s -960 228156 480 228396 4 io_in[18]
port 9 nsew signal input
rlabel metal2 s 204598 619520 204710 620960 6 io_in[19]
port 10 nsew signal input
rlabel metal2 s 42310 -960 42422 480 8 io_in[1]
port 11 nsew signal input
rlabel metal2 s 149950 619520 150062 620960 6 io_in[20]
port 12 nsew signal input
rlabel metal2 s 174238 619520 174350 620960 6 io_in[21]
port 13 nsew signal input
rlabel metal3 s -960 62508 480 62748 4 io_in[22]
port 14 nsew signal input
rlabel metal3 s -960 169948 480 170188 4 io_in[23]
port 15 nsew signal input
rlabel metal3 s 499520 447388 500960 447628 6 io_in[24]
port 16 nsew signal input
rlabel metal2 s 50038 619520 50150 620960 6 io_in[25]
port 17 nsew signal input
rlabel metal2 s 325670 619520 325782 620960 6 io_in[26]
port 18 nsew signal input
rlabel metal2 s 159150 619520 159262 620960 6 io_in[27]
port 19 nsew signal input
rlabel metal3 s -960 26604 480 26844 4 io_in[28]
port 20 nsew signal input
rlabel metal2 s 243974 619520 244086 620960 6 io_in[29]
port 21 nsew signal input
rlabel metal3 s -960 555100 480 555340 4 io_in[2]
port 22 nsew signal input
rlabel metal2 s 196686 -960 196798 480 8 io_in[30]
port 23 nsew signal input
rlabel metal3 s -960 196876 480 197116 4 io_in[31]
port 24 nsew signal input
rlabel metal2 s 349958 619520 350070 620960 6 io_in[32]
port 25 nsew signal input
rlabel metal2 s 304510 619520 304622 620960 6 io_in[33]
port 26 nsew signal input
rlabel metal2 s 139278 -960 139390 480 8 io_in[34]
port 27 nsew signal input
rlabel metal3 s 499520 393532 500960 393772 6 io_in[35]
port 28 nsew signal input
rlabel metal3 s -960 232508 480 232748 4 io_in[36]
port 29 nsew signal input
rlabel metal2 s 427054 -960 427166 480 8 io_in[37]
port 30 nsew signal input
rlabel metal3 s -960 237132 480 237372 4 io_in[3]
port 31 nsew signal input
rlabel metal2 s 474158 619520 474270 620960 6 io_in[4]
port 32 nsew signal input
rlabel metal3 s 499520 30956 500960 31196 6 io_in[5]
port 33 nsew signal input
rlabel metal3 s 499520 344300 500960 344540 6 io_in[6]
port 34 nsew signal input
rlabel metal3 s -960 375852 480 376092 4 io_in[7]
port 35 nsew signal input
rlabel metal2 s 255934 619520 256046 620960 6 io_in[8]
port 36 nsew signal input
rlabel metal3 s -960 438684 480 438924 4 io_in[9]
port 37 nsew signal input
rlabel metal3 s 499520 187628 500960 187868 6 io_oeb[0]
port 38 nsew signal tristate
rlabel metal3 s 499520 174300 500960 174540 6 io_oeb[10]
port 39 nsew signal tristate
rlabel metal2 s 310582 619520 310694 620960 6 io_oeb[11]
port 40 nsew signal tristate
rlabel metal2 s 195398 619520 195510 620960 6 io_oeb[12]
port 41 nsew signal tristate
rlabel metal2 s 342230 -960 342342 480 8 io_oeb[13]
port 42 nsew signal tristate
rlabel metal2 s 113702 619520 113814 620960 6 io_oeb[14]
port 43 nsew signal tristate
rlabel metal3 s 499520 191980 500960 192220 6 io_oeb[15]
port 44 nsew signal tristate
rlabel metal2 s 314814 -960 314926 480 8 io_oeb[16]
port 45 nsew signal tristate
rlabel metal2 s 34950 619520 35062 620960 6 io_oeb[17]
port 46 nsew signal tristate
rlabel metal2 s 43966 619520 44078 620960 6 io_oeb[18]
port 47 nsew signal tristate
rlabel metal3 s -960 205852 480 206092 4 io_oeb[19]
port 48 nsew signal tristate
rlabel metal2 s 311870 -960 311982 480 8 io_oeb[1]
port 49 nsew signal tristate
rlabel metal2 s 116646 619520 116758 620960 6 io_oeb[20]
port 50 nsew signal tristate
rlabel metal2 s 352902 619520 353014 620960 6 io_oeb[21]
port 51 nsew signal tristate
rlabel metal3 s -960 120716 480 120956 4 io_oeb[22]
port 52 nsew signal tristate
rlabel metal3 s 499520 223532 500960 223772 6 io_oeb[23]
port 53 nsew signal tristate
rlabel metal3 s 499520 613036 500960 613276 6 io_oeb[24]
port 54 nsew signal tristate
rlabel metal3 s -960 528172 480 528412 4 io_oeb[25]
port 55 nsew signal tristate
rlabel metal2 s 86470 619520 86582 620960 6 io_oeb[26]
port 56 nsew signal tristate
rlabel metal3 s -960 8652 480 8892 4 io_oeb[27]
port 57 nsew signal tristate
rlabel metal2 s 316654 619520 316766 620960 6 io_oeb[28]
port 58 nsew signal tristate
rlabel metal3 s 499520 442764 500960 443004 6 io_oeb[29]
port 59 nsew signal tristate
rlabel metal3 s 499520 527900 500960 528140 6 io_oeb[2]
port 60 nsew signal tristate
rlabel metal2 s 287582 -960 287694 480 8 io_oeb[30]
port 61 nsew signal tristate
rlabel metal3 s -960 595356 480 595596 4 io_oeb[31]
port 62 nsew signal tristate
rlabel metal2 s 92358 619520 92470 620960 6 io_oeb[32]
port 63 nsew signal tristate
rlabel metal2 s 52982 619520 53094 620960 6 io_oeb[33]
port 64 nsew signal tristate
rlabel metal2 s 119774 619520 119886 620960 6 io_oeb[34]
port 65 nsew signal tristate
rlabel metal3 s -960 366876 480 367116 4 io_oeb[35]
port 66 nsew signal tristate
rlabel metal2 s 205886 -960 205998 480 8 io_oeb[36]
port 67 nsew signal tristate
rlabel metal3 s -960 496892 480 497132 4 io_oeb[37]
port 68 nsew signal tristate
rlabel metal2 s 389334 619520 389446 620960 6 io_oeb[3]
port 69 nsew signal tristate
rlabel metal2 s 233118 -960 233230 480 8 io_oeb[4]
port 70 nsew signal tristate
rlabel metal3 s -960 183276 480 183516 4 io_oeb[5]
port 71 nsew signal tristate
rlabel metal2 s 367990 619520 368102 620960 6 io_oeb[6]
port 72 nsew signal tristate
rlabel metal2 s 483174 619520 483286 620960 6 io_oeb[7]
port 73 nsew signal tristate
rlabel metal3 s -960 478940 480 479180 4 io_oeb[8]
port 74 nsew signal tristate
rlabel metal2 s 80398 619520 80510 620960 6 io_oeb[9]
port 75 nsew signal tristate
rlabel metal2 s 28878 619520 28990 620960 6 io_out[0]
port 76 nsew signal tristate
rlabel metal2 s 471030 619520 471142 620960 6 io_out[10]
port 77 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_out[11]
port 78 nsew signal tristate
rlabel metal3 s 499520 572780 500960 573020 6 io_out[12]
port 79 nsew signal tristate
rlabel metal3 s -960 219180 480 219420 4 io_out[13]
port 80 nsew signal tristate
rlabel metal2 s 60526 -960 60638 480 8 io_out[14]
port 81 nsew signal tristate
rlabel metal3 s 499520 469692 500960 469932 6 io_out[15]
port 82 nsew signal tristate
rlabel metal3 s 499520 102492 500960 102732 6 io_out[16]
port 83 nsew signal tristate
rlabel metal3 s 499520 384556 500960 384796 6 io_out[17]
port 84 nsew signal tristate
rlabel metal3 s 499520 550204 500960 550444 6 io_out[18]
port 85 nsew signal tristate
rlabel metal3 s 499520 474316 500960 474556 6 io_out[19]
port 86 nsew signal tristate
rlabel metal2 s 54454 -960 54566 480 8 io_out[1]
port 87 nsew signal tristate
rlabel metal2 s 354190 -960 354302 480 8 io_out[20]
port 88 nsew signal tristate
rlabel metal2 s 22806 619520 22918 620960 6 io_out[21]
port 89 nsew signal tristate
rlabel metal2 s 439014 -960 439126 480 8 io_out[22]
port 90 nsew signal tristate
rlabel metal2 s 257406 -960 257518 480 8 io_out[23]
port 91 nsew signal tristate
rlabel metal3 s 499520 21980 500960 22220 6 io_out[24]
port 92 nsew signal tristate
rlabel metal3 s -960 460988 480 461228 4 io_out[25]
port 93 nsew signal tristate
rlabel metal2 s 125846 619520 125958 620960 6 io_out[26]
port 94 nsew signal tristate
rlabel metal2 s 463302 -960 463414 480 8 io_out[27]
port 95 nsew signal tristate
rlabel metal3 s 499520 321996 500960 322236 6 io_out[28]
port 96 nsew signal tristate
rlabel metal2 s 108918 -960 109030 480 8 io_out[29]
port 97 nsew signal tristate
rlabel metal2 s 480230 619520 480342 620960 6 io_out[2]
port 98 nsew signal tristate
rlabel metal2 s 145350 -960 145462 480 8 io_out[30]
port 99 nsew signal tristate
rlabel metal3 s 499520 541228 500960 541468 6 io_out[31]
port 100 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 io_out[32]
port 101 nsew signal tristate
rlabel metal3 s 499520 456364 500960 456604 6 io_out[33]
port 102 nsew signal tristate
rlabel metal2 s 495318 619520 495430 620960 6 io_out[34]
port 103 nsew signal tristate
rlabel metal3 s 499520 402508 500960 402748 6 io_out[35]
port 104 nsew signal tristate
rlabel metal2 s 122718 619520 122830 620960 6 io_out[36]
port 105 nsew signal tristate
rlabel metal2 s 414910 -960 415022 480 8 io_out[37]
port 106 nsew signal tristate
rlabel metal3 s -960 331244 480 331484 4 io_out[3]
port 107 nsew signal tristate
rlabel metal3 s 499520 13004 500960 13244 6 io_out[4]
port 108 nsew signal tristate
rlabel metal3 s 499520 366604 500960 366844 6 io_out[5]
port 109 nsew signal tristate
rlabel metal2 s 268078 619520 268190 620960 6 io_out[6]
port 110 nsew signal tristate
rlabel metal3 s -960 156620 480 156860 4 io_out[7]
port 111 nsew signal tristate
rlabel metal2 s 222630 619520 222742 620960 6 io_out[8]
port 112 nsew signal tristate
rlabel metal2 s 25750 619520 25862 620960 6 io_out[9]
port 113 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 irq[0]
port 114 nsew signal tristate
rlabel metal3 s 499520 218908 500960 219148 6 irq[1]
port 115 nsew signal tristate
rlabel metal2 s 401478 619520 401590 620960 6 irq[2]
port 116 nsew signal tristate
rlabel metal3 s 499520 290716 500960 290956 6 la_data_in[0]
port 117 nsew signal input
rlabel metal3 s 499520 138396 500960 138636 6 la_data_in[100]
port 118 nsew signal input
rlabel metal2 s 237902 619520 238014 620960 6 la_data_in[101]
port 119 nsew signal input
rlabel metal2 s 107630 619520 107742 620960 6 la_data_in[102]
port 120 nsew signal input
rlabel metal3 s 499520 563804 500960 564044 6 la_data_in[103]
port 121 nsew signal input
rlabel metal3 s -960 510220 480 510460 4 la_data_in[104]
port 122 nsew signal input
rlabel metal3 s 499520 371228 500960 371468 6 la_data_in[105]
port 123 nsew signal input
rlabel metal3 s 499520 17356 500960 17596 6 la_data_in[106]
port 124 nsew signal input
rlabel metal2 s 286294 619520 286406 620960 6 la_data_in[107]
port 125 nsew signal input
rlabel metal3 s 499520 125068 500960 125308 6 la_data_in[108]
port 126 nsew signal input
rlabel metal2 s 365046 619520 365158 620960 6 la_data_in[109]
port 127 nsew signal input
rlabel metal3 s -960 523548 480 523788 4 la_data_in[10]
port 128 nsew signal input
rlabel metal2 s 15078 -960 15190 480 8 la_data_in[110]
port 129 nsew signal input
rlabel metal3 s 499520 375580 500960 375820 6 la_data_in[111]
port 130 nsew signal input
rlabel metal3 s -960 532524 480 532764 4 la_data_in[112]
port 131 nsew signal input
rlabel metal3 s 499520 53260 500960 53500 6 la_data_in[113]
port 132 nsew signal input
rlabel metal2 s 377190 619520 377302 620960 6 la_data_in[114]
port 133 nsew signal input
rlabel metal2 s 112046 -960 112158 480 8 la_data_in[115]
port 134 nsew signal input
rlabel metal2 s 202758 -960 202870 480 8 la_data_in[116]
port 135 nsew signal input
rlabel metal2 s 219686 619520 219798 620960 6 la_data_in[117]
port 136 nsew signal input
rlabel metal2 s 407366 619520 407478 620960 6 la_data_in[118]
port 137 nsew signal input
rlabel metal3 s 499520 353276 500960 353516 6 la_data_in[119]
port 138 nsew signal input
rlabel metal3 s -960 487916 480 488156 4 la_data_in[11]
port 139 nsew signal input
rlabel metal2 s 346830 619520 346942 620960 6 la_data_in[120]
port 140 nsew signal input
rlabel metal2 s 448214 -960 448326 480 8 la_data_in[121]
port 141 nsew signal input
rlabel metal2 s 56110 619520 56222 620960 6 la_data_in[122]
port 142 nsew signal input
rlabel metal2 s 469374 -960 469486 480 8 la_data_in[123]
port 143 nsew signal input
rlabel metal2 s 74326 619520 74438 620960 6 la_data_in[124]
port 144 nsew signal input
rlabel metal3 s -960 174300 480 174540 4 la_data_in[125]
port 145 nsew signal input
rlabel metal2 s 351246 -960 351358 480 8 la_data_in[126]
port 146 nsew signal input
rlabel metal3 s -960 362524 480 362764 4 la_data_in[127]
port 147 nsew signal input
rlabel metal3 s -960 304316 480 304556 4 la_data_in[12]
port 148 nsew signal input
rlabel metal2 s 408838 -960 408950 480 8 la_data_in[13]
port 149 nsew signal input
rlabel metal3 s 499520 433788 500960 434028 6 la_data_in[14]
port 150 nsew signal input
rlabel metal3 s -960 107388 480 107628 4 la_data_in[15]
port 151 nsew signal input
rlabel metal3 s 499520 232508 500960 232748 6 la_data_in[16]
port 152 nsew signal input
rlabel metal3 s -960 277388 480 277628 4 la_data_in[17]
port 153 nsew signal input
rlabel metal3 s 499520 514572 500960 514812 6 la_data_in[18]
port 154 nsew signal input
rlabel metal2 s 386206 619520 386318 620960 6 la_data_in[19]
port 155 nsew signal input
rlabel metal2 s 114990 -960 115102 480 8 la_data_in[1]
port 156 nsew signal input
rlabel metal2 s 41022 619520 41134 620960 6 la_data_in[20]
port 157 nsew signal input
rlabel metal3 s -960 22252 480 22492 4 la_data_in[21]
port 158 nsew signal input
rlabel metal2 s 305798 -960 305910 480 8 la_data_in[22]
port 159 nsew signal input
rlabel metal3 s 499520 304044 500960 304284 6 la_data_in[23]
port 160 nsew signal input
rlabel metal3 s 499520 80188 500960 80428 6 la_data_in[24]
port 161 nsew signal input
rlabel metal3 s -960 447660 480 447900 4 la_data_in[25]
port 162 nsew signal input
rlabel metal3 s 499520 487644 500960 487884 6 la_data_in[26]
port 163 nsew signal input
rlabel metal3 s -960 49180 480 49420 4 la_data_in[27]
port 164 nsew signal input
rlabel metal3 s 499520 348924 500960 349164 6 la_data_in[28]
port 165 nsew signal input
rlabel metal2 s 330086 -960 330198 480 8 la_data_in[29]
port 166 nsew signal input
rlabel metal2 s 366334 -960 366446 480 8 la_data_in[2]
port 167 nsew signal input
rlabel metal2 s 432942 -960 433054 480 8 la_data_in[30]
port 168 nsew signal input
rlabel metal2 s 201470 619520 201582 620960 6 la_data_in[31]
port 169 nsew signal input
rlabel metal2 s 336158 -960 336270 480 8 la_data_in[32]
port 170 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[33]
port 171 nsew signal input
rlabel metal2 s 246918 619520 247030 620960 6 la_data_in[34]
port 172 nsew signal input
rlabel metal3 s -960 564076 480 564316 4 la_data_in[35]
port 173 nsew signal input
rlabel metal2 s 398350 619520 398462 620960 6 la_data_in[36]
port 174 nsew signal input
rlabel metal2 s 486118 619520 486230 620960 6 la_data_in[37]
port 175 nsew signal input
rlabel metal3 s 499520 241484 500960 241724 6 la_data_in[38]
port 176 nsew signal input
rlabel metal2 s 9006 -960 9118 480 8 la_data_in[39]
port 177 nsew signal input
rlabel metal3 s -960 348924 480 349164 4 la_data_in[3]
port 178 nsew signal input
rlabel metal2 s 93830 -960 93942 480 8 la_data_in[40]
port 179 nsew signal input
rlabel metal2 s 121062 -960 121174 480 8 la_data_in[41]
port 180 nsew signal input
rlabel metal3 s 499520 254812 500960 255052 6 la_data_in[42]
port 181 nsew signal input
rlabel metal3 s 499520 465340 500960 465580 6 la_data_in[43]
port 182 nsew signal input
rlabel metal2 s 186382 619520 186494 620960 6 la_data_in[44]
port 183 nsew signal input
rlabel metal3 s -960 116092 480 116332 4 la_data_in[45]
port 184 nsew signal input
rlabel metal3 s -960 371500 480 371740 4 la_data_in[46]
port 185 nsew signal input
rlabel metal2 s 308926 -960 309038 480 8 la_data_in[47]
port 186 nsew signal input
rlabel metal2 s 362102 619520 362214 620960 6 la_data_in[48]
port 187 nsew signal input
rlabel metal2 s 90702 -960 90814 480 8 la_data_in[49]
port 188 nsew signal input
rlabel metal2 s 160438 -960 160550 480 8 la_data_in[4]
port 189 nsew signal input
rlabel metal3 s -960 13276 480 13516 4 la_data_in[50]
port 190 nsew signal input
rlabel metal2 s 37894 619520 38006 620960 6 la_data_in[51]
port 191 nsew signal input
rlabel metal2 s 477102 619520 477214 620960 6 la_data_in[52]
port 192 nsew signal input
rlabel metal3 s 499520 75564 500960 75804 6 la_data_in[53]
port 193 nsew signal input
rlabel metal2 s 57398 -960 57510 480 8 la_data_in[54]
port 194 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[55]
port 195 nsew signal input
rlabel metal2 s 2934 -960 3046 480 8 la_data_in[56]
port 196 nsew signal input
rlabel metal2 s 345174 -960 345286 480 8 la_data_in[57]
port 197 nsew signal input
rlabel metal2 s 419510 619520 419622 620960 6 la_data_in[58]
port 198 nsew signal input
rlabel metal2 s 402766 -960 402878 480 8 la_data_in[59]
port 199 nsew signal input
rlabel metal3 s -960 286364 480 286604 4 la_data_in[5]
port 200 nsew signal input
rlabel metal2 s 68254 619520 68366 620960 6 la_data_in[60]
port 201 nsew signal input
rlabel metal2 s 96774 -960 96886 480 8 la_data_in[61]
port 202 nsew signal input
rlabel metal3 s 499520 111468 500960 111708 6 la_data_in[62]
port 203 nsew signal input
rlabel metal3 s -960 380476 480 380716 4 la_data_in[63]
port 204 nsew signal input
rlabel metal3 s 499520 581756 500960 581996 6 la_data_in[64]
port 205 nsew signal input
rlabel metal2 s 399638 -960 399750 480 8 la_data_in[65]
port 206 nsew signal input
rlabel metal2 s 10662 619520 10774 620960 6 la_data_in[66]
port 207 nsew signal input
rlabel metal2 s 225758 619520 225870 620960 6 la_data_in[67]
port 208 nsew signal input
rlabel metal3 s -960 165596 480 165836 4 la_data_in[68]
port 209 nsew signal input
rlabel metal3 s 499520 438412 500960 438652 6 la_data_in[69]
port 210 nsew signal input
rlabel metal3 s 499520 214556 500960 214796 6 la_data_in[6]
port 211 nsew signal input
rlabel metal3 s 499520 116092 500960 116332 6 la_data_in[70]
port 212 nsew signal input
rlabel metal3 s 499520 71212 500960 71452 6 la_data_in[71]
port 213 nsew signal input
rlabel metal2 s 147006 619520 147118 620960 6 la_data_in[72]
port 214 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_data_in[73]
port 215 nsew signal input
rlabel metal2 s 227046 -960 227158 480 8 la_data_in[74]
port 216 nsew signal input
rlabel metal2 s 181598 -960 181710 480 8 la_data_in[75]
port 217 nsew signal input
rlabel metal2 s 224102 -960 224214 480 8 la_data_in[76]
port 218 nsew signal input
rlabel metal3 s 499520 380204 500960 380444 6 la_data_in[77]
port 219 nsew signal input
rlabel metal3 s 499520 483020 500960 483260 6 la_data_in[78]
port 220 nsew signal input
rlabel metal3 s 499520 133772 500960 134012 6 la_data_in[79]
port 221 nsew signal input
rlabel metal3 s 499520 156348 500960 156588 6 la_data_in[7]
port 222 nsew signal input
rlabel metal2 s 378478 -960 378590 480 8 la_data_in[80]
port 223 nsew signal input
rlabel metal3 s 499520 160700 500960 160940 6 la_data_in[81]
port 224 nsew signal input
rlabel metal3 s -960 299692 480 299932 4 la_data_in[82]
port 225 nsew signal input
rlabel metal2 s 422638 619520 422750 620960 6 la_data_in[83]
port 226 nsew signal input
rlabel metal3 s -960 4300 480 4540 4 la_data_in[84]
port 227 nsew signal input
rlabel metal2 s 216558 619520 216670 620960 6 la_data_in[85]
port 228 nsew signal input
rlabel metal3 s 499520 424812 500960 425052 6 la_data_in[86]
port 229 nsew signal input
rlabel metal3 s -960 340220 480 340460 4 la_data_in[87]
port 230 nsew signal input
rlabel metal3 s -960 411756 480 411996 4 la_data_in[88]
port 231 nsew signal input
rlabel metal2 s 192454 619520 192566 620960 6 la_data_in[89]
port 232 nsew signal input
rlabel metal2 s 140934 619520 141046 620960 6 la_data_in[8]
port 233 nsew signal input
rlabel metal2 s 301382 619520 301494 620960 6 la_data_in[90]
port 234 nsew signal input
rlabel metal2 s 47094 619520 47206 620960 6 la_data_in[91]
port 235 nsew signal input
rlabel metal2 s 472318 -960 472430 480 8 la_data_in[92]
port 236 nsew signal input
rlabel metal2 s 163382 -960 163494 480 8 la_data_in[93]
port 237 nsew signal input
rlabel metal2 s 184726 -960 184838 480 8 la_data_in[94]
port 238 nsew signal input
rlabel metal3 s 499520 4028 500960 4268 6 la_data_in[95]
port 239 nsew signal input
rlabel metal3 s -960 241484 480 241724 4 la_data_in[96]
port 240 nsew signal input
rlabel metal3 s -960 590732 480 590972 4 la_data_in[97]
port 241 nsew signal input
rlabel metal3 s 499520 263788 500960 264028 6 la_data_in[98]
port 242 nsew signal input
rlabel metal3 s -960 456636 480 456876 4 la_data_in[99]
port 243 nsew signal input
rlabel metal2 s 81686 -960 81798 480 8 la_data_in[9]
port 244 nsew signal input
rlabel metal3 s -960 425084 480 425324 4 la_data_out[0]
port 245 nsew signal tristate
rlabel metal2 s 464958 619520 465070 620960 6 la_data_out[100]
port 246 nsew signal tristate
rlabel metal3 s -960 586380 480 586620 4 la_data_out[101]
port 247 nsew signal tristate
rlabel metal3 s -960 57884 480 58124 4 la_data_out[102]
port 248 nsew signal tristate
rlabel metal3 s 499520 196604 500960 196844 6 la_data_out[103]
port 249 nsew signal tristate
rlabel metal3 s 499520 313020 500960 313260 6 la_data_out[104]
port 250 nsew signal tristate
rlabel metal3 s -960 214828 480 215068 4 la_data_out[105]
port 251 nsew signal tristate
rlabel metal2 s 137806 619520 137918 620960 6 la_data_out[106]
port 252 nsew signal tristate
rlabel metal2 s 302854 -960 302966 480 8 la_data_out[107]
port 253 nsew signal tristate
rlabel metal3 s -960 537148 480 537388 4 la_data_out[108]
port 254 nsew signal tristate
rlabel metal2 s 274150 619520 274262 620960 6 la_data_out[109]
port 255 nsew signal tristate
rlabel metal2 s 313526 619520 313638 620960 6 la_data_out[10]
port 256 nsew signal tristate
rlabel metal2 s 72670 -960 72782 480 8 la_data_out[110]
port 257 nsew signal tristate
rlabel metal2 s 374062 619520 374174 620960 6 la_data_out[111]
port 258 nsew signal tristate
rlabel metal2 s 455942 619520 456054 620960 6 la_data_out[112]
port 259 nsew signal tristate
rlabel metal3 s -960 53532 480 53772 4 la_data_out[113]
port 260 nsew signal tristate
rlabel metal2 s 228702 619520 228814 620960 6 la_data_out[114]
port 261 nsew signal tristate
rlabel metal3 s 499520 536876 500960 537116 6 la_data_out[115]
port 262 nsew signal tristate
rlabel metal3 s 499520 98140 500960 98380 6 la_data_out[116]
port 263 nsew signal tristate
rlabel metal3 s -960 160972 480 161212 4 la_data_out[117]
port 264 nsew signal tristate
rlabel metal2 s 175526 -960 175638 480 8 la_data_out[118]
port 265 nsew signal tristate
rlabel metal3 s -960 246108 480 246348 4 la_data_out[119]
port 266 nsew signal tristate
rlabel metal2 s 263478 -960 263590 480 8 la_data_out[11]
port 267 nsew signal tristate
rlabel metal2 s 478390 -960 478502 480 8 la_data_out[120]
port 268 nsew signal tristate
rlabel metal2 s 110574 619520 110686 620960 6 la_data_out[121]
port 269 nsew signal tristate
rlabel metal2 s 462014 619520 462126 620960 6 la_data_out[122]
port 270 nsew signal tristate
rlabel metal3 s -960 541500 480 541740 4 la_data_out[123]
port 271 nsew signal tristate
rlabel metal3 s -960 223804 480 224044 4 la_data_out[124]
port 272 nsew signal tristate
rlabel metal2 s 420982 -960 421094 480 8 la_data_out[125]
port 273 nsew signal tristate
rlabel metal2 s 266422 -960 266534 480 8 la_data_out[126]
port 274 nsew signal tristate
rlabel metal3 s -960 407132 480 407372 4 la_data_out[127]
port 275 nsew signal tristate
rlabel metal3 s 499520 545852 500960 546092 6 la_data_out[12]
port 276 nsew signal tristate
rlabel metal3 s 499520 250188 500960 250428 6 la_data_out[13]
port 277 nsew signal tristate
rlabel metal3 s -960 264060 480 264300 4 la_data_out[14]
port 278 nsew signal tristate
rlabel metal3 s 499520 281740 500960 281980 6 la_data_out[15]
port 279 nsew signal tristate
rlabel metal2 s 454286 -960 454398 480 8 la_data_out[16]
port 280 nsew signal tristate
rlabel metal2 s 71198 619520 71310 620960 6 la_data_out[17]
port 281 nsew signal tristate
rlabel metal3 s 499520 62236 500960 62476 6 la_data_out[18]
port 282 nsew signal tristate
rlabel metal3 s -960 434060 480 434300 4 la_data_out[19]
port 283 nsew signal tristate
rlabel metal2 s 65126 619520 65238 620960 6 la_data_out[1]
port 284 nsew signal tristate
rlabel metal3 s 499520 599436 500960 599676 6 la_data_out[20]
port 285 nsew signal tristate
rlabel metal3 s -960 138668 480 138908 4 la_data_out[21]
port 286 nsew signal tristate
rlabel metal2 s 337814 619520 337926 620960 6 la_data_out[22]
port 287 nsew signal tristate
rlabel metal3 s 499520 200956 500960 201196 6 la_data_out[23]
port 288 nsew signal tristate
rlabel metal2 s 211958 -960 212070 480 8 la_data_out[24]
port 289 nsew signal tristate
rlabel metal2 s 292366 619520 292478 620960 6 la_data_out[25]
port 290 nsew signal tristate
rlabel metal3 s -960 134044 480 134284 4 la_data_out[26]
port 291 nsew signal tristate
rlabel metal3 s 499520 259164 500960 259404 6 la_data_out[27]
port 292 nsew signal tristate
rlabel metal2 s 69542 -960 69654 480 8 la_data_out[28]
port 293 nsew signal tristate
rlabel metal2 s 4590 619520 4702 620960 6 la_data_out[29]
port 294 nsew signal tristate
rlabel metal3 s 499520 44284 500960 44524 6 la_data_out[2]
port 295 nsew signal tristate
rlabel metal2 s 214902 -960 215014 480 8 la_data_out[30]
port 296 nsew signal tristate
rlabel metal3 s -960 201228 480 201468 4 la_data_out[31]
port 297 nsew signal tristate
rlabel metal2 s 131734 619520 131846 620960 6 la_data_out[32]
port 298 nsew signal tristate
rlabel metal2 s 298438 619520 298550 620960 6 la_data_out[33]
port 299 nsew signal tristate
rlabel metal2 s 445086 -960 445198 480 8 la_data_out[34]
port 300 nsew signal tristate
rlabel metal2 s 443798 619520 443910 620960 6 la_data_out[35]
port 301 nsew signal tristate
rlabel metal3 s -960 505868 480 506108 4 la_data_out[36]
port 302 nsew signal tristate
rlabel metal3 s -960 322268 480 322508 4 la_data_out[37]
port 303 nsew signal tristate
rlabel metal2 s 404422 619520 404534 620960 6 la_data_out[38]
port 304 nsew signal tristate
rlabel metal3 s 499520 129420 500960 129660 6 la_data_out[39]
port 305 nsew signal tristate
rlabel metal2 s 210486 619520 210598 620960 6 la_data_out[3]
port 306 nsew signal tristate
rlabel metal3 s -960 429708 480 429948 4 la_data_out[40]
port 307 nsew signal tristate
rlabel metal2 s 260350 -960 260462 480 8 la_data_out[41]
port 308 nsew signal tristate
rlabel metal2 s 177182 619520 177294 620960 6 la_data_out[42]
port 309 nsew signal tristate
rlabel metal2 s 162094 619520 162206 620960 6 la_data_out[43]
port 310 nsew signal tristate
rlabel metal2 s 387678 -960 387790 480 8 la_data_out[44]
port 311 nsew signal tristate
rlabel metal2 s 475446 -960 475558 480 8 la_data_out[45]
port 312 nsew signal tristate
rlabel metal2 s 492190 619520 492302 620960 6 la_data_out[46]
port 313 nsew signal tristate
rlabel metal2 s 198526 619520 198638 620960 6 la_data_out[47]
port 314 nsew signal tristate
rlabel metal3 s -960 80460 480 80700 4 la_data_out[48]
port 315 nsew signal tristate
rlabel metal2 s 33294 -960 33406 480 8 la_data_out[49]
port 316 nsew signal tristate
rlabel metal3 s -960 317644 480 317884 4 la_data_out[4]
port 317 nsew signal tristate
rlabel metal3 s -960 384828 480 385068 4 la_data_out[50]
port 318 nsew signal tristate
rlabel metal2 s 142222 -960 142334 480 8 la_data_out[51]
port 319 nsew signal tristate
rlabel metal3 s -960 514844 480 515084 4 la_data_out[52]
port 320 nsew signal tristate
rlabel metal3 s 499520 286092 500960 286332 6 la_data_out[53]
port 321 nsew signal tristate
rlabel metal3 s -960 416108 480 416348 4 la_data_out[54]
port 322 nsew signal tristate
rlabel metal3 s 499520 268140 500960 268380 6 la_data_out[55]
port 323 nsew signal tristate
rlabel metal3 s -960 35580 480 35820 4 la_data_out[56]
port 324 nsew signal tristate
rlabel metal2 s 242134 -960 242246 480 8 la_data_out[57]
port 325 nsew signal tristate
rlabel metal2 s 468086 619520 468198 620960 6 la_data_out[58]
port 326 nsew signal tristate
rlabel metal2 s 392278 619520 392390 620960 6 la_data_out[59]
port 327 nsew signal tristate
rlabel metal2 s 259062 619520 259174 620960 6 la_data_out[5]
port 328 nsew signal tristate
rlabel metal2 s 63470 -960 63582 480 8 la_data_out[60]
port 329 nsew signal tristate
rlabel metal2 s 363390 -960 363502 480 8 la_data_out[61]
port 330 nsew signal tristate
rlabel metal3 s -960 577404 480 577644 4 la_data_out[62]
port 331 nsew signal tristate
rlabel metal3 s 499520 308396 500960 308636 6 la_data_out[63]
port 332 nsew signal tristate
rlabel metal3 s 499520 93516 500960 93756 6 la_data_out[64]
port 333 nsew signal tristate
rlabel metal3 s 499520 35308 500960 35548 6 la_data_out[65]
port 334 nsew signal tristate
rlabel metal2 s 220974 -960 221086 480 8 la_data_out[66]
port 335 nsew signal tristate
rlabel metal2 s 326958 -960 327070 480 8 la_data_out[67]
port 336 nsew signal tristate
rlabel metal2 s 169454 -960 169566 480 8 la_data_out[68]
port 337 nsew signal tristate
rlabel metal2 s 452814 619520 452926 620960 6 la_data_out[69]
port 338 nsew signal tristate
rlabel metal2 s 251334 -960 251446 480 8 la_data_out[6]
port 339 nsew signal tristate
rlabel metal2 s 213614 619520 213726 620960 6 la_data_out[70]
port 340 nsew signal tristate
rlabel metal2 s 13606 619520 13718 620960 6 la_data_out[71]
port 341 nsew signal tristate
rlabel metal2 s 124006 -960 124118 480 8 la_data_out[72]
port 342 nsew signal tristate
rlabel metal2 s 265134 619520 265246 620960 6 la_data_out[73]
port 343 nsew signal tristate
rlabel metal2 s 230174 -960 230286 480 8 la_data_out[74]
port 344 nsew signal tristate
rlabel metal3 s 499520 8652 500960 8892 6 la_data_out[75]
port 345 nsew signal tristate
rlabel metal2 s 436070 -960 436182 480 8 la_data_out[76]
port 346 nsew signal tristate
rlabel metal3 s 499520 89164 500960 89404 6 la_data_out[77]
port 347 nsew signal tristate
rlabel metal3 s 499520 57884 500960 58124 6 la_data_out[78]
port 348 nsew signal tristate
rlabel metal2 s 172582 -960 172694 480 8 la_data_out[79]
port 349 nsew signal tristate
rlabel metal2 s 1646 619520 1758 620960 6 la_data_out[7]
port 350 nsew signal tristate
rlabel metal3 s -960 84812 480 85052 4 la_data_out[80]
port 351 nsew signal tristate
rlabel metal2 s 134862 619520 134974 620960 6 la_data_out[81]
port 352 nsew signal tristate
rlabel metal2 s 375534 -960 375646 480 8 la_data_out[82]
port 353 nsew signal tristate
rlabel metal2 s 101558 619520 101670 620960 6 la_data_out[83]
port 354 nsew signal tristate
rlabel metal3 s -960 125068 480 125308 4 la_data_out[84]
port 355 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[85]
port 356 nsew signal tristate
rlabel metal3 s 499520 295068 500960 295308 6 la_data_out[86]
port 357 nsew signal tristate
rlabel metal2 s 289238 619520 289350 620960 6 la_data_out[87]
port 358 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[88]
port 359 nsew signal tristate
rlabel metal2 s 277278 619520 277390 620960 6 la_data_out[89]
port 360 nsew signal tristate
rlabel metal2 s 280222 619520 280334 620960 6 la_data_out[8]
port 361 nsew signal tristate
rlabel metal2 s 348302 -960 348414 480 8 la_data_out[90]
port 362 nsew signal tristate
rlabel metal2 s 390622 -960 390734 480 8 la_data_out[91]
port 363 nsew signal tristate
rlabel metal2 s 428710 619520 428822 620960 6 la_data_out[92]
port 364 nsew signal tristate
rlabel metal2 s 183254 619520 183366 620960 6 la_data_out[93]
port 365 nsew signal tristate
rlabel metal2 s 231830 619520 231942 620960 6 la_data_out[94]
port 366 nsew signal tristate
rlabel metal2 s 360262 -960 360374 480 8 la_data_out[95]
port 367 nsew signal tristate
rlabel metal2 s 77270 619520 77382 620960 6 la_data_out[96]
port 368 nsew signal tristate
rlabel metal3 s -960 255084 480 255324 4 la_data_out[97]
port 369 nsew signal tristate
rlabel metal2 s 416566 619520 416678 620960 6 la_data_out[98]
port 370 nsew signal tristate
rlabel metal2 s 466430 -960 466542 480 8 la_data_out[99]
port 371 nsew signal tristate
rlabel metal2 s 208830 -960 208942 480 8 la_data_out[9]
port 372 nsew signal tristate
rlabel metal2 s 245262 -960 245374 480 8 la_oenb[0]
port 373 nsew signal input
rlabel metal3 s 499520 608412 500960 608652 6 la_oenb[100]
port 374 nsew signal input
rlabel metal3 s -960 568428 480 568668 4 la_oenb[101]
port 375 nsew signal input
rlabel metal2 s 425582 619520 425694 620960 6 la_oenb[102]
port 376 nsew signal input
rlabel metal2 s 117934 -960 118046 480 8 la_oenb[103]
port 377 nsew signal input
rlabel metal3 s 499520 335324 500960 335564 6 la_oenb[104]
port 378 nsew signal input
rlabel metal2 s 249862 619520 249974 620960 6 la_oenb[105]
port 379 nsew signal input
rlabel metal2 s 489246 619520 489358 620960 6 la_oenb[106]
port 380 nsew signal input
rlabel metal3 s 499520 326348 500960 326588 6 la_oenb[107]
port 381 nsew signal input
rlabel metal2 s 340758 619520 340870 620960 6 la_oenb[108]
port 382 nsew signal input
rlabel metal2 s 395406 619520 395518 620960 6 la_oenb[109]
port 383 nsew signal input
rlabel metal2 s 187670 -960 187782 480 8 la_oenb[10]
port 384 nsew signal input
rlabel metal3 s 499520 460716 500960 460956 6 la_oenb[110]
port 385 nsew signal input
rlabel metal2 s 339102 -960 339214 480 8 la_oenb[111]
port 386 nsew signal input
rlabel metal3 s -960 353548 480 353788 4 la_oenb[112]
port 387 nsew signal input
rlabel metal2 s 87758 -960 87870 480 8 la_oenb[113]
port 388 nsew signal input
rlabel metal2 s 307454 619520 307566 620960 6 la_oenb[114]
port 389 nsew signal input
rlabel metal2 s 269550 -960 269662 480 8 la_oenb[115]
port 390 nsew signal input
rlabel metal2 s 239190 -960 239302 480 8 la_oenb[116]
port 391 nsew signal input
rlabel metal3 s 499520 586108 500960 586348 6 la_oenb[117]
port 392 nsew signal input
rlabel metal3 s 499520 209932 500960 210172 6 la_oenb[118]
port 393 nsew signal input
rlabel metal3 s -960 326620 480 326860 4 la_oenb[119]
port 394 nsew signal input
rlabel metal3 s 499520 330972 500960 331212 6 la_oenb[11]
port 395 nsew signal input
rlabel metal2 s 296782 -960 296894 480 8 la_oenb[120]
port 396 nsew signal input
rlabel metal2 s 166510 -960 166622 480 8 la_oenb[121]
port 397 nsew signal input
rlabel metal3 s -960 492268 480 492508 4 la_oenb[122]
port 398 nsew signal input
rlabel metal3 s 499520 505596 500960 505836 6 la_oenb[123]
port 399 nsew signal input
rlabel metal3 s -960 393804 480 394044 4 la_oenb[124]
port 400 nsew signal input
rlabel metal3 s -960 465340 480 465580 4 la_oenb[125]
port 401 nsew signal input
rlabel metal2 s 381606 -960 381718 480 8 la_oenb[126]
port 402 nsew signal input
rlabel metal3 s 499520 120444 500960 120684 6 la_oenb[127]
port 403 nsew signal input
rlabel metal3 s 499520 411484 500960 411724 6 la_oenb[12]
port 404 nsew signal input
rlabel metal3 s -960 111740 480 111980 4 la_oenb[13]
port 405 nsew signal input
rlabel metal3 s -960 93788 480 94028 4 la_oenb[14]
port 406 nsew signal input
rlabel metal2 s 248206 -960 248318 480 8 la_oenb[15]
port 407 nsew signal input
rlabel metal2 s 133206 -960 133318 480 8 la_oenb[16]
port 408 nsew signal input
rlabel metal3 s 499520 66860 500960 67100 6 la_oenb[17]
port 409 nsew signal input
rlabel metal2 s 30166 -960 30278 480 8 la_oenb[18]
port 410 nsew signal input
rlabel metal2 s 136150 -960 136262 480 8 la_oenb[19]
port 411 nsew signal input
rlabel metal3 s 499520 48908 500960 49148 6 la_oenb[1]
port 412 nsew signal input
rlabel metal3 s 499520 577132 500960 577372 6 la_oenb[20]
port 413 nsew signal input
rlabel metal3 s 499520 227884 500960 228124 6 la_oenb[21]
port 414 nsew signal input
rlabel metal2 s 48382 -960 48494 480 8 la_oenb[22]
port 415 nsew signal input
rlabel metal3 s -960 210204 480 210444 4 la_oenb[23]
port 416 nsew signal input
rlabel metal2 s 324014 -960 324126 480 8 la_oenb[24]
port 417 nsew signal input
rlabel metal2 s 440854 619520 440966 620960 6 la_oenb[25]
port 418 nsew signal input
rlabel metal2 s 299726 -960 299838 480 8 la_oenb[26]
port 419 nsew signal input
rlabel metal3 s 499520 317372 500960 317612 6 la_oenb[27]
port 420 nsew signal input
rlabel metal2 s 498262 619520 498374 620960 6 la_oenb[28]
port 421 nsew signal input
rlabel metal2 s 446742 619520 446854 620960 6 la_oenb[29]
port 422 nsew signal input
rlabel metal3 s -960 31228 480 31468 4 la_oenb[2]
port 423 nsew signal input
rlabel metal3 s -960 313292 480 313532 4 la_oenb[30]
port 424 nsew signal input
rlabel metal2 s 168166 619520 168278 620960 6 la_oenb[31]
port 425 nsew signal input
rlabel metal2 s 154366 -960 154478 480 8 la_oenb[32]
port 426 nsew signal input
rlabel metal2 s 89414 619520 89526 620960 6 la_oenb[33]
port 427 nsew signal input
rlabel metal3 s 499520 165324 500960 165564 6 la_oenb[34]
port 428 nsew signal input
rlabel metal3 s 499520 339948 500960 340188 6 la_oenb[35]
port 429 nsew signal input
rlabel metal3 s -960 89436 480 89676 4 la_oenb[36]
port 430 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oenb[37]
port 431 nsew signal input
rlabel metal3 s 499520 496620 500960 496860 6 la_oenb[38]
port 432 nsew signal input
rlabel metal3 s -960 452012 480 452252 4 la_oenb[39]
port 433 nsew signal input
rlabel metal2 s 458886 619520 458998 620960 6 la_oenb[3]
port 434 nsew signal input
rlabel metal3 s -960 581756 480 581996 4 la_oenb[40]
port 435 nsew signal input
rlabel metal2 s 429998 -960 430110 480 8 la_oenb[41]
port 436 nsew signal input
rlabel metal2 s 59054 619520 59166 620960 6 la_oenb[42]
port 437 nsew signal input
rlabel metal3 s -960 573052 480 573292 4 la_oenb[43]
port 438 nsew signal input
rlabel metal2 s 493662 -960 493774 480 8 la_oenb[44]
port 439 nsew signal input
rlabel metal2 s 84630 -960 84742 480 8 la_oenb[45]
port 440 nsew signal input
rlabel metal2 s 127134 -960 127246 480 8 la_oenb[46]
port 441 nsew signal input
rlabel metal2 s 442142 -960 442254 480 8 la_oenb[47]
port 442 nsew signal input
rlabel metal3 s 499520 151724 500960 151964 6 la_oenb[48]
port 443 nsew signal input
rlabel metal3 s 499520 500972 500960 501212 6 la_oenb[49]
port 444 nsew signal input
rlabel metal3 s -960 469964 480 470204 4 la_oenb[4]
port 445 nsew signal input
rlabel metal2 s 252990 619520 253102 620960 6 la_oenb[50]
port 446 nsew signal input
rlabel metal2 s 180310 619520 180422 620960 6 la_oenb[51]
port 447 nsew signal input
rlabel metal3 s -960 335596 480 335836 4 la_oenb[52]
port 448 nsew signal input
rlabel metal3 s 499520 568156 500960 568396 6 la_oenb[53]
port 449 nsew signal input
rlabel metal3 s -960 501244 480 501484 4 la_oenb[54]
port 450 nsew signal input
rlabel metal2 s 153078 619520 153190 620960 6 la_oenb[55]
port 451 nsew signal input
rlabel metal3 s -960 98412 480 98652 4 la_oenb[56]
port 452 nsew signal input
rlabel metal3 s 499520 491996 500960 492236 6 la_oenb[57]
port 453 nsew signal input
rlabel metal2 s 358974 619520 359086 620960 6 la_oenb[58]
port 454 nsew signal input
rlabel metal2 s 7718 619520 7830 620960 6 la_oenb[59]
port 455 nsew signal input
rlabel metal2 s 410494 619520 410606 620960 6 la_oenb[5]
port 456 nsew signal input
rlabel metal2 s 434782 619520 434894 620960 6 la_oenb[60]
port 457 nsew signal input
rlabel metal2 s 437726 619520 437838 620960 6 la_oenb[61]
port 458 nsew signal input
rlabel metal2 s 275438 -960 275550 480 8 la_oenb[62]
port 459 nsew signal input
rlabel metal2 s 283350 619520 283462 620960 6 la_oenb[63]
port 460 nsew signal input
rlabel metal2 s 18022 -960 18134 480 8 la_oenb[64]
port 461 nsew signal input
rlabel metal2 s 5878 -960 5990 480 8 la_oenb[65]
port 462 nsew signal input
rlabel metal2 s 411782 -960 411894 480 8 la_oenb[66]
port 463 nsew signal input
rlabel metal3 s -960 282012 480 282252 4 la_oenb[67]
port 464 nsew signal input
rlabel metal3 s 499520 84540 500960 84780 6 la_oenb[68]
port 465 nsew signal input
rlabel metal3 s -960 357900 480 358140 4 la_oenb[69]
port 466 nsew signal input
rlabel metal3 s -960 474316 480 474556 4 la_oenb[6]
port 467 nsew signal input
rlabel metal2 s 19678 619520 19790 620960 6 la_oenb[70]
port 468 nsew signal input
rlabel metal3 s -960 295340 480 295580 4 la_oenb[71]
port 469 nsew signal input
rlabel metal3 s -960 250460 480 250700 4 la_oenb[72]
port 470 nsew signal input
rlabel metal3 s -960 192252 480 192492 4 la_oenb[73]
port 471 nsew signal input
rlabel metal2 s 271206 619520 271318 620960 6 la_oenb[74]
port 472 nsew signal input
rlabel metal2 s 423926 -960 424038 480 8 la_oenb[75]
port 473 nsew signal input
rlabel metal2 s 199814 -960 199926 480 8 la_oenb[76]
port 474 nsew signal input
rlabel metal3 s -960 550476 480 550716 4 la_oenb[77]
port 475 nsew signal input
rlabel metal3 s 499520 416108 500960 416348 6 la_oenb[78]
port 476 nsew signal input
rlabel metal3 s 499520 559180 500960 559420 6 la_oenb[79]
port 477 nsew signal input
rlabel metal3 s -960 398428 480 398668 4 la_oenb[7]
port 478 nsew signal input
rlabel metal3 s -960 483292 480 483532 4 la_oenb[80]
port 479 nsew signal input
rlabel metal3 s 499520 26332 500960 26572 6 la_oenb[81]
port 480 nsew signal input
rlabel metal3 s 499520 523548 500960 523788 6 la_oenb[82]
port 481 nsew signal input
rlabel metal2 s 207542 619520 207654 620960 6 la_oenb[83]
port 482 nsew signal input
rlabel metal3 s 499520 429436 500960 429676 6 la_oenb[84]
port 483 nsew signal input
rlabel metal2 s 396694 -960 396806 480 8 la_oenb[85]
port 484 nsew signal input
rlabel metal3 s -960 344572 480 344812 4 la_oenb[86]
port 485 nsew signal input
rlabel metal3 s 499520 107116 500960 107356 6 la_oenb[87]
port 486 nsew signal input
rlabel metal2 s 171110 619520 171222 620960 6 la_oenb[88]
port 487 nsew signal input
rlabel metal2 s 481518 -960 481630 480 8 la_oenb[89]
port 488 nsew signal input
rlabel metal3 s -960 613308 480 613548 4 la_oenb[8]
port 489 nsew signal input
rlabel metal2 s 66598 -960 66710 480 8 la_oenb[90]
port 490 nsew signal input
rlabel metal3 s -960 259436 480 259676 4 la_oenb[91]
port 491 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_oenb[92]
port 492 nsew signal input
rlabel metal3 s 499520 518924 500960 519164 6 la_oenb[93]
port 493 nsew signal input
rlabel metal2 s 130078 -960 130190 480 8 la_oenb[94]
port 494 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_oenb[95]
port 495 nsew signal input
rlabel metal2 s 31822 619520 31934 620960 6 la_oenb[96]
port 496 nsew signal input
rlabel metal2 s 322726 619520 322838 620960 6 la_oenb[97]
port 497 nsew signal input
rlabel metal3 s -960 102764 480 103004 4 la_oenb[98]
port 498 nsew signal input
rlabel metal2 s 16734 619520 16846 620960 6 la_oenb[99]
port 499 nsew signal input
rlabel metal2 s 62182 619520 62294 620960 6 la_oenb[9]
port 500 nsew signal input
rlabel metal3 s 499520 147372 500960 147612 6 wb_clk_i
port 501 nsew signal input
rlabel metal3 s -960 604332 480 604572 4 wb_rst_i
port 502 nsew signal input
rlabel metal3 s -960 187900 480 188140 4 wbs_ack_o
port 503 nsew signal tristate
rlabel metal2 s 234774 619520 234886 620960 6 wbs_adr_i[0]
port 504 nsew signal input
rlabel metal2 s 128790 619520 128902 620960 6 wbs_adr_i[10]
port 505 nsew signal input
rlabel metal3 s -960 519196 480 519436 4 wbs_adr_i[11]
port 506 nsew signal input
rlabel metal2 s 45254 -960 45366 480 8 wbs_adr_i[12]
port 507 nsew signal input
rlabel metal3 s -960 402780 480 403020 4 wbs_adr_i[13]
port 508 nsew signal input
rlabel metal3 s 499520 554828 500960 555068 6 wbs_adr_i[14]
port 509 nsew signal input
rlabel metal3 s 499520 509948 500960 510188 6 wbs_adr_i[15]
port 510 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 wbs_adr_i[16]
port 511 nsew signal input
rlabel metal3 s -960 44556 480 44796 4 wbs_adr_i[17]
port 512 nsew signal input
rlabel metal3 s 499520 236860 500960 237100 6 wbs_adr_i[18]
port 513 nsew signal input
rlabel metal2 s 484462 -960 484574 480 8 wbs_adr_i[19]
port 514 nsew signal input
rlabel metal2 s 240846 619520 240958 620960 6 wbs_adr_i[1]
port 515 nsew signal input
rlabel metal2 s 383262 619520 383374 620960 6 wbs_adr_i[20]
port 516 nsew signal input
rlabel metal2 s 284638 -960 284750 480 8 wbs_adr_i[21]
port 517 nsew signal input
rlabel metal2 s 405710 -960 405822 480 8 wbs_adr_i[22]
port 518 nsew signal input
rlabel metal3 s 499520 169676 500960 169916 6 wbs_adr_i[23]
port 519 nsew signal input
rlabel metal3 s -960 599708 480 599948 4 wbs_adr_i[24]
port 520 nsew signal input
rlabel metal2 s 272494 -960 272606 480 8 wbs_adr_i[25]
port 521 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[26]
port 522 nsew signal input
rlabel metal2 s 98430 619520 98542 620960 6 wbs_adr_i[27]
port 523 nsew signal input
rlabel metal3 s 499520 420460 500960 420700 6 wbs_adr_i[28]
port 524 nsew signal input
rlabel metal2 s 449870 619520 449982 620960 6 wbs_adr_i[29]
port 525 nsew signal input
rlabel metal2 s 193742 -960 193854 480 8 wbs_adr_i[2]
port 526 nsew signal input
rlabel metal2 s 328614 619520 328726 620960 6 wbs_adr_i[30]
port 527 nsew signal input
rlabel metal3 s 499520 299692 500960 299932 6 wbs_adr_i[31]
port 528 nsew signal input
rlabel metal2 s 384550 -960 384662 480 8 wbs_adr_i[3]
port 529 nsew signal input
rlabel metal2 s 319598 619520 319710 620960 6 wbs_adr_i[4]
port 530 nsew signal input
rlabel metal2 s 369462 -960 369574 480 8 wbs_adr_i[5]
port 531 nsew signal input
rlabel metal2 s 157310 -960 157422 480 8 wbs_adr_i[6]
port 532 nsew signal input
rlabel metal2 s 24094 -960 24206 480 8 wbs_adr_i[7]
port 533 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 wbs_adr_i[8]
port 534 nsew signal input
rlabel metal3 s 499520 183276 500960 183516 6 wbs_adr_i[9]
port 535 nsew signal input
rlabel metal2 s 104502 619520 104614 620960 6 wbs_cyc_i
port 536 nsew signal input
rlabel metal3 s 499520 617388 500960 617628 6 wbs_dat_i[0]
port 537 nsew signal input
rlabel metal3 s -960 389452 480 389692 4 wbs_dat_i[10]
port 538 nsew signal input
rlabel metal3 s -960 443036 480 443276 4 wbs_dat_i[11]
port 539 nsew signal input
rlabel metal3 s -960 66860 480 67100 4 wbs_dat_i[12]
port 540 nsew signal input
rlabel metal2 s 21150 -960 21262 480 8 wbs_dat_i[13]
port 541 nsew signal input
rlabel metal2 s 105974 -960 106086 480 8 wbs_dat_i[14]
port 542 nsew signal input
rlabel metal3 s 499520 357900 500960 358140 6 wbs_dat_i[15]
port 543 nsew signal input
rlabel metal2 s 278566 -960 278678 480 8 wbs_dat_i[16]
port 544 nsew signal input
rlabel metal2 s 295310 619520 295422 620960 6 wbs_dat_i[17]
port 545 nsew signal input
rlabel metal2 s 413438 619520 413550 620960 6 wbs_dat_i[18]
port 546 nsew signal input
rlabel metal3 s -960 608684 480 608924 4 wbs_dat_i[19]
port 547 nsew signal input
rlabel metal2 s 75614 -960 75726 480 8 wbs_dat_i[1]
port 548 nsew signal input
rlabel metal3 s 499520 407132 500960 407372 6 wbs_dat_i[20]
port 549 nsew signal input
rlabel metal2 s 431654 619520 431766 620960 6 wbs_dat_i[21]
port 550 nsew signal input
rlabel metal3 s -960 290716 480 290956 4 wbs_dat_i[22]
port 551 nsew signal input
rlabel metal3 s 499520 532524 500960 532764 6 wbs_dat_i[23]
port 552 nsew signal input
rlabel metal3 s 499520 205580 500960 205820 6 wbs_dat_i[24]
port 553 nsew signal input
rlabel metal3 s -960 17628 480 17868 4 wbs_dat_i[25]
port 554 nsew signal input
rlabel metal2 s 380134 619520 380246 620960 6 wbs_dat_i[26]
port 555 nsew signal input
rlabel metal2 s 95486 619520 95598 620960 6 wbs_dat_i[27]
port 556 nsew signal input
rlabel metal2 s 151422 -960 151534 480 8 wbs_dat_i[28]
port 557 nsew signal input
rlabel metal3 s 499520 398156 500960 398396 6 wbs_dat_i[29]
port 558 nsew signal input
rlabel metal2 s 393566 -960 393678 480 8 wbs_dat_i[2]
port 559 nsew signal input
rlabel metal3 s 499520 178652 500960 178892 6 wbs_dat_i[30]
port 560 nsew signal input
rlabel metal3 s -960 268412 480 268652 4 wbs_dat_i[31]
port 561 nsew signal input
rlabel metal2 s 496606 -960 496718 480 8 wbs_dat_i[3]
port 562 nsew signal input
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_i[4]
port 563 nsew signal input
rlabel metal2 s 236062 -960 236174 480 8 wbs_dat_i[5]
port 564 nsew signal input
rlabel metal3 s 499520 272764 500960 273004 6 wbs_dat_i[6]
port 565 nsew signal input
rlabel metal2 s 371118 619520 371230 620960 6 wbs_dat_i[7]
port 566 nsew signal input
rlabel metal3 s 499520 595084 500960 595324 6 wbs_dat_i[8]
port 567 nsew signal input
rlabel metal2 s 499734 -960 499846 480 8 wbs_dat_i[9]
port 568 nsew signal input
rlabel metal2 s 39182 -960 39294 480 8 wbs_dat_o[0]
port 569 nsew signal tristate
rlabel metal3 s 499520 362252 500960 362492 6 wbs_dat_o[10]
port 570 nsew signal tristate
rlabel metal2 s 11950 -960 12062 480 8 wbs_dat_o[11]
port 571 nsew signal tristate
rlabel metal3 s 499520 604060 500960 604300 6 wbs_dat_o[12]
port 572 nsew signal tristate
rlabel metal2 s 356030 619520 356142 620960 6 wbs_dat_o[13]
port 573 nsew signal tristate
rlabel metal3 s 499520 39932 500960 40172 6 wbs_dat_o[14]
port 574 nsew signal tristate
rlabel metal3 s -960 75836 480 76076 4 wbs_dat_o[15]
port 575 nsew signal tristate
rlabel metal3 s -960 129692 480 129932 4 wbs_dat_o[16]
port 576 nsew signal tristate
rlabel metal3 s -960 151996 480 152236 4 wbs_dat_o[17]
port 577 nsew signal tristate
rlabel metal2 s 317942 -960 318054 480 8 wbs_dat_o[18]
port 578 nsew signal tristate
rlabel metal2 s -10 -960 102 480 8 wbs_dat_o[19]
port 579 nsew signal tristate
rlabel metal2 s 372406 -960 372518 480 8 wbs_dat_o[1]
port 580 nsew signal tristate
rlabel metal3 s -960 273036 480 273276 4 wbs_dat_o[20]
port 581 nsew signal tristate
rlabel metal3 s -960 546124 480 546364 4 wbs_dat_o[21]
port 582 nsew signal tristate
rlabel metal2 s 143878 619520 143990 620960 6 wbs_dat_o[22]
port 583 nsew signal tristate
rlabel metal3 s -960 178924 480 179164 4 wbs_dat_o[23]
port 584 nsew signal tristate
rlabel metal2 s 99902 -960 100014 480 8 wbs_dat_o[24]
port 585 nsew signal tristate
rlabel metal2 s 36238 -960 36350 480 8 wbs_dat_o[25]
port 586 nsew signal tristate
rlabel metal2 s 262006 619520 262118 620960 6 wbs_dat_o[26]
port 587 nsew signal tristate
rlabel metal2 s 156022 619520 156134 620960 6 wbs_dat_o[27]
port 588 nsew signal tristate
rlabel metal2 s 254278 -960 254390 480 8 wbs_dat_o[28]
port 589 nsew signal tristate
rlabel metal2 s 343886 619520 343998 620960 6 wbs_dat_o[29]
port 590 nsew signal tristate
rlabel metal3 s 499520 142748 500960 142988 6 wbs_dat_o[2]
port 591 nsew signal tristate
rlabel metal3 s -960 420732 480 420972 4 wbs_dat_o[30]
port 592 nsew signal tristate
rlabel metal3 s 499520 478668 500960 478908 6 wbs_dat_o[31]
port 593 nsew signal tristate
rlabel metal2 s 102846 -960 102958 480 8 wbs_dat_o[3]
port 594 nsew signal tristate
rlabel metal2 s 178654 -960 178766 480 8 wbs_dat_o[4]
port 595 nsew signal tristate
rlabel metal3 s -960 40204 480 40444 4 wbs_dat_o[5]
port 596 nsew signal tristate
rlabel metal3 s 499520 451740 500960 451980 6 wbs_dat_o[6]
port 597 nsew signal tristate
rlabel metal2 s 281510 -960 281622 480 8 wbs_dat_o[7]
port 598 nsew signal tristate
rlabel metal2 s 334686 619520 334798 620960 6 wbs_dat_o[8]
port 599 nsew signal tristate
rlabel metal2 s 331742 619520 331854 620960 6 wbs_dat_o[9]
port 600 nsew signal tristate
rlabel metal3 s -960 617660 480 617900 4 wbs_sel_i[0]
port 601 nsew signal input
rlabel metal2 s 83342 619520 83454 620960 6 wbs_sel_i[1]
port 602 nsew signal input
rlabel metal2 s 333030 -960 333142 480 8 wbs_sel_i[2]
port 603 nsew signal input
rlabel metal3 s -960 143020 480 143260 4 wbs_sel_i[3]
port 604 nsew signal input
rlabel metal3 s -960 559452 480 559692 4 wbs_stb_i
port 605 nsew signal input
rlabel metal3 s 499520 277116 500960 277356 6 wbs_we_i
port 606 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 500000 620000
<< end >>
